module vop_decoder (
    input                   clk,
    input                   reset,
    input                   stall,
    input [1:0][9:0]        opcodes,
    output reg [1:0][3:0]   vops
);

always_comb begin // lane 1
    vops[0] = 9; // default to NOP
    case (opcodes[0])
        46: vops[0] = 0; // DADDU
        67: vops[0] = 0; // DSRAV
        47: vops[0] = 0; // DSUB
        89: vops[0] = 0; // DMULT_LO
        92: vops[0] = 0; // DMULTU_HI
        86: vops[0] = 0; // MULT_HI
        73: vops[0] = 0; // DDIV_HI
        68: vops[0] = 0; // DIV_LO
        71: vops[0] = 0; // DIVU_HI
        36: vops[0] = 0; // ADDU
        54: vops[0] = 0; // SLLV
        41: vops[0] = 0; // SLTU
        39: vops[0] = 0; // OR
        361: vops[0] = 0; // MOVN_1
        360: vops[0] = 0; // MOVN_0
        74: vops[0] = 0; // DDIVU_LO
        48: vops[0] = 0; // DSUBU
        88: vops[0] = 0; // MULTU_HI
        40: vops[0] = 0; // SLT
        52: vops[0] = 0; // ROTRV
        43: vops[0] = 0; // SUBU
        37: vops[0] = 0; // AND
        61: vops[0] = 0; // DSLLV
        38: vops[0] = 0; // NOR
        84: vops[0] = 0; // MUL
        91: vops[0] = 0; // DMULTU_LO
        64: vops[0] = 0; // DSRLV
        90: vops[0] = 0; // DMULT_HI
        85: vops[0] = 0; // MULT_LO
        368: vops[0] = 0; // MOVZ_1
        367: vops[0] = 0; // MOVZ_0
        70: vops[0] = 0; // DIVU_LO
        69: vops[0] = 0; // DIV_HI
        72: vops[0] = 0; // DDIV_LO
        58: vops[0] = 0; // SRLV
        75: vops[0] = 0; // DDIVU_HI
        56: vops[0] = 0; // SRAV
        87: vops[0] = 0; // MULTU_LO
        44: vops[0] = 0; // XOR
        45: vops[0] = 0; // DADD
        137: vops[0] = 1; // EXT
        139: vops[0] = 1; // DEXT
        62: vops[0] = 1; // DSRL
        65: vops[0] = 1; // DSRA
        30: vops[0] = 1; // SLTI
        63: vops[0] = 1; // DSRL32
        53: vops[0] = 1; // SLL
        59: vops[0] = 1; // DSLL
        60: vops[0] = 1; // DSLL32
        27: vops[0] = 1; // ANDI
        55: vops[0] = 1; // SRA
        57: vops[0] = 1; // SRL
        34: vops[0] = 1; // DADDIU
        32: vops[0] = 1; // XORI
        31: vops[0] = 1; // SLTIU
        29: vops[0] = 1; // ORI
        51: vops[0] = 1; // ROTR
        66: vops[0] = 1; // DSRA32
        26: vops[0] = 1; // ADDIU
        141: vops[0] = 1; // DEXTU
        140: vops[0] = 1; // DEXTM
        81: vops[0] = 2; // MSUBU
        80: vops[0] = 2; // MSUB
        76: vops[0] = 2; // MADD
        77: vops[0] = 2; // MADDU
        119: vops[0] = 3; // SYSCALL
        118: vops[0] = 3; // BREAK
        122: vops[0] = 4; // TGEU
        120: vops[0] = 4; // TEQ
        123: vops[0] = 4; // TLT
        124: vops[0] = 4; // TLTU
        121: vops[0] = 4; // TGE
        125: vops[0] = 4; // TNE
        127: vops[0] = 5; // TGEI
        126: vops[0] = 5; // TEQI
        128: vops[0] = 5; // TGEIU
        131: vops[0] = 5; // TNEI
        129: vops[0] = 5; // TLTI
        130: vops[0] = 5; // TLTIU
        136: vops[0] = 6; // EHB
        25: vops[0] = 7; // ADDI
        33: vops[0] = 7; // DADDI
        78: vops[0] = 8; // MFHI
        147: vops[0] = 8; // WSBH
        83: vops[0] = 8; // MTLO
        145: vops[0] = 8; // SEB
        50: vops[0] = 8; // CLZ
        146: vops[0] = 8; // SEH
        79: vops[0] = 8; // MFLO
        49: vops[0] = 8; // CLO
        82: vops[0] = 8; // MTHI
        116: vops[0] = 9; // SYNC
        134: vops[0] = 9; // NOP
        135: vops[0] = 9; // SSNOP
        138: vops[0] = 10; // INS
        142: vops[0] = 10; // DINS
        144: vops[0] = 10; // DINSU
        143: vops[0] = 10; // DINSM
        153: vops[0] = 11; // RDHWR
        28: vops[0] = 11; // LUI
        42: vops[0] = 12; // SUB
        35: vops[0] = 12; // ADD
        117: vops[0] = 13; // SYNCI
        1: vops[0] = 0; // LBU
        3: vops[0] = 0; // LHU
        20: vops[0] = 0; // LLD
        5: vops[0] = 0; // LWU
        9: vops[0] = 0; // LD
        0: vops[0] = 0; // LB
        19: vops[0] = 0; // LL
        2: vops[0] = 0; // LH
        4: vops[0] = 0; // LW
        14: vops[0] = 1; // LDR
        13: vops[0] = 1; // LDL
        12: vops[0] = 1; // LWR
        11: vops[0] = 1; // LWL
        133: vops[0] = 2; // PREFX
        132: vops[0] = 2; // PREF
        22: vops[0] = 0; // SC_1
        24: vops[0] = 0; // SCD_1
        21: vops[0] = 1; // SC_0
        23: vops[0] = 1; // SCD_0
        8: vops[0] = 1; // SW
        7: vops[0] = 1; // SH
        6: vops[0] = 1; // SB
        10: vops[0] = 1; // SD
        15: vops[0] = 1; // SWL
        16: vops[0] = 1; // SWR
        17: vops[0] = 1; // SDL
        18: vops[0] = 1; // SDR
        98: vops[0] = 0; // JR
        99: vops[0] = 0; // JR_HB
        115: vops[0] = 1; // BNEL
        101: vops[0] = 1; // BNE
        100: vops[0] = 1; // BEQ
        108: vops[0] = 1; // BEQL
        106: vops[0] = 2; // BLTZ
        111: vops[0] = 2; // BGTZL
        114: vops[0] = 2; // BLTZL
        105: vops[0] = 2; // BLEZ
        110: vops[0] = 2; // BGEZL
        112: vops[0] = 2; // BLEZL
        102: vops[0] = 2; // BGEZ
        104: vops[0] = 2; // BGTZ
        97: vops[0] = 3; // JALR_HB
        96: vops[0] = 3; // JALR
        113: vops[0] = 4; // BLTZALL
        109: vops[0] = 4; // BGEZALL
        103: vops[0] = 4; // BGEZAL
        107: vops[0] = 4; // BLTZAL
        93: vops[0] = 5; // J
        95: vops[0] = 6; // JALX
        94: vops[0] = 6; // JAL
    endcase // opcodes[0]
end

always_comb begin // lane 2
    vops[1] = 9; // default to NOP
    case (opcodes[1])
        46: vops[1] = 0; // DADDU
        67: vops[1] = 0; // DSRAV
        47: vops[1] = 0; // DSUB
        89: vops[1] = 0; // DMULT_LO
        92: vops[1] = 0; // DMULTU_HI
        86: vops[1] = 0; // MULT_HI
        73: vops[1] = 0; // DDIV_HI
        68: vops[1] = 0; // DIV_LO
        71: vops[1] = 0; // DIVU_HI
        36: vops[1] = 0; // ADDU
        54: vops[1] = 0; // SLLV
        41: vops[1] = 0; // SLTU
        39: vops[1] = 0; // OR
        361: vops[1] = 0; // MOVN_1
        360: vops[1] = 0; // MOVN_0
        74: vops[1] = 0; // DDIVU_LO
        48: vops[1] = 0; // DSUBU
        88: vops[1] = 0; // MULTU_HI
        40: vops[1] = 0; // SLT
        52: vops[1] = 0; // ROTRV
        43: vops[1] = 0; // SUBU
        37: vops[1] = 0; // AND
        61: vops[1] = 0; // DSLLV
        38: vops[1] = 0; // NOR
        84: vops[1] = 0; // MUL
        91: vops[1] = 0; // DMULTU_LO
        64: vops[1] = 0; // DSRLV
        90: vops[1] = 0; // DMULT_HI
        85: vops[1] = 0; // MULT_LO
        368: vops[1] = 0; // MOVZ_1
        367: vops[1] = 0; // MOVZ_0
        70: vops[1] = 0; // DIVU_LO
        69: vops[1] = 0; // DIV_HI
        72: vops[1] = 0; // DDIV_LO
        58: vops[1] = 0; // SRLV
        75: vops[1] = 0; // DDIVU_HI
        56: vops[1] = 0; // SRAV
        87: vops[1] = 0; // MULTU_LO
        44: vops[1] = 0; // XOR
        45: vops[1] = 0; // DADD
        137: vops[1] = 1; // EXT
        139: vops[1] = 1; // DEXT
        62: vops[1] = 1; // DSRL
        65: vops[1] = 1; // DSRA
        30: vops[1] = 1; // SLTI
        63: vops[1] = 1; // DSRL32
        53: vops[1] = 1; // SLL
        59: vops[1] = 1; // DSLL
        60: vops[1] = 1; // DSLL32
        27: vops[1] = 1; // ANDI
        55: vops[1] = 1; // SRA
        57: vops[1] = 1; // SRL
        34: vops[1] = 1; // DADDIU
        32: vops[1] = 1; // XORI
        31: vops[1] = 1; // SLTIU
        29: vops[1] = 1; // ORI
        51: vops[1] = 1; // ROTR
        66: vops[1] = 1; // DSRA32
        26: vops[1] = 1; // ADDIU
        141: vops[1] = 1; // DEXTU
        140: vops[1] = 1; // DEXTM
        81: vops[1] = 2; // MSUBU
        80: vops[1] = 2; // MSUB
        76: vops[1] = 2; // MADD
        77: vops[1] = 2; // MADDU
        119: vops[1] = 3; // SYSCALL
        118: vops[1] = 3; // BREAK
        122: vops[1] = 4; // TGEU
        120: vops[1] = 4; // TEQ
        123: vops[1] = 4; // TLT
        124: vops[1] = 4; // TLTU
        121: vops[1] = 4; // TGE
        125: vops[1] = 4; // TNE
        127: vops[1] = 5; // TGEI
        126: vops[1] = 5; // TEQI
        128: vops[1] = 5; // TGEIU
        131: vops[1] = 5; // TNEI
        129: vops[1] = 5; // TLTI
        130: vops[1] = 5; // TLTIU
        136: vops[1] = 6; // EHB
        25: vops[1] = 7; // ADDI
        33: vops[1] = 7; // DADDI
        78: vops[1] = 8; // MFHI
        147: vops[1] = 8; // WSBH
        83: vops[1] = 8; // MTLO
        145: vops[1] = 8; // SEB
        50: vops[1] = 8; // CLZ
        146: vops[1] = 8; // SEH
        79: vops[1] = 8; // MFLO
        49: vops[1] = 8; // CLO
        82: vops[1] = 8; // MTHI
        116: vops[1] = 9; // SYNC
        134: vops[1] = 9; // NOP
        135: vops[1] = 9; // SSNOP
        138: vops[1] = 10; // INS
        142: vops[1] = 10; // DINS
        144: vops[1] = 10; // DINSU
        143: vops[1] = 10; // DINSM
        153: vops[1] = 11; // RDHWR
        28: vops[1] = 11; // LUI
        42: vops[1] = 12; // SUB
        35: vops[1] = 12; // ADD
        117: vops[1] = 13; // SYNCI
        1: vops[1] = 0; // LBU
        3: vops[1] = 0; // LHU
        20: vops[1] = 0; // LLD
        5: vops[1] = 0; // LWU
        9: vops[1] = 0; // LD
        0: vops[1] = 0; // LB
        19: vops[1] = 0; // LL
        2: vops[1] = 0; // LH
        4: vops[1] = 0; // LW
        14: vops[1] = 1; // LDR
        13: vops[1] = 1; // LDL
        12: vops[1] = 1; // LWR
        11: vops[1] = 1; // LWL
        133: vops[1] = 2; // PREFX
        132: vops[1] = 2; // PREF
        22: vops[1] = 0; // SC_1
        24: vops[1] = 0; // SCD_1
        21: vops[1] = 1; // SC_0
        23: vops[1] = 1; // SCD_0
        8: vops[1] = 1; // SW
        7: vops[1] = 1; // SH
        6: vops[1] = 1; // SB
        10: vops[1] = 1; // SD
        15: vops[1] = 1; // SWL
        16: vops[1] = 1; // SWR
        17: vops[1] = 1; // SDL
        18: vops[1] = 1; // SDR
        98: vops[1] = 0; // JR
        99: vops[1] = 0; // JR_HB
        115: vops[1] = 1; // BNEL
        101: vops[1] = 1; // BNE
        100: vops[1] = 1; // BEQ
        108: vops[1] = 1; // BEQL
        106: vops[1] = 2; // BLTZ
        111: vops[1] = 2; // BGTZL
        114: vops[1] = 2; // BLTZL
        105: vops[1] = 2; // BLEZ
        110: vops[1] = 2; // BGEZL
        112: vops[1] = 2; // BLEZL
        102: vops[1] = 2; // BGEZ
        104: vops[1] = 2; // BGTZ
        97: vops[1] = 3; // JALR_HB
        96: vops[1] = 3; // JALR
        113: vops[1] = 4; // BLTZALL
        109: vops[1] = 4; // BGEZALL
        103: vops[1] = 4; // BGEZAL
        107: vops[1] = 4; // BLTZAL
        93: vops[1] = 5; // J
        95: vops[1] = 6; // JALX
        94: vops[1] = 6; // JAL
    endcase // opcodes[1]
end

endmodule
