module ecc_checker_10(data_in, checker_in, parity_in);

input      [ 501:0] data_in;
output reg [  8:0] checker_in;
output reg         parity_in;

always @(*) begin
    checker_in[0] = data_in[501] ^ data_in[500] ^ data_in[498] ^ data_in[497] ^ data_in[495] ^ data_in[493] ^ data_in[491] ^ data_in[490] ^ data_in[488] ^ data_in[486] ^ data_in[484] ^ data_in[482] ^ data_in[480] ^ data_in[478] ^ data_in[476] ^ data_in[475] ^ data_in[473] ^ data_in[471] ^ data_in[469] ^ data_in[467] ^ data_in[465] ^ data_in[463] ^ data_in[461] ^ data_in[459] ^ data_in[457] ^ data_in[455] ^ data_in[453] ^ data_in[451] ^ data_in[449] ^ data_in[447] ^ data_in[445] ^ data_in[444] ^ data_in[442] ^ data_in[440] ^ data_in[438] ^ data_in[436] ^ data_in[434] ^ data_in[432] ^ data_in[430] ^ data_in[428] ^ data_in[426] ^ data_in[424] ^ data_in[422] ^ data_in[420] ^ data_in[418] ^ data_in[416] ^ data_in[414] ^ data_in[412] ^ data_in[410] ^ data_in[408] ^ data_in[406] ^ data_in[404] ^ data_in[402] ^ data_in[400] ^ data_in[398] ^ data_in[396] ^ data_in[394] ^ data_in[392] ^ data_in[390] ^ data_in[388] ^ data_in[386] ^ data_in[384] ^ data_in[382] ^ data_in[381] ^ data_in[379] ^ data_in[377] ^ data_in[375] ^ data_in[373] ^ data_in[371] ^ data_in[369] ^ data_in[367] ^ data_in[365] ^ data_in[363] ^ data_in[361] ^ data_in[359] ^ data_in[357] ^ data_in[355] ^ data_in[353] ^ data_in[351] ^ data_in[349] ^ data_in[347] ^ data_in[345] ^ data_in[343] ^ data_in[341] ^ data_in[339] ^ data_in[337] ^ data_in[335] ^ data_in[333] ^ data_in[331] ^ data_in[329] ^ data_in[327] ^ data_in[325] ^ data_in[323] ^ data_in[321] ^ data_in[319] ^ data_in[317] ^ data_in[315] ^ data_in[313] ^ data_in[311] ^ data_in[309] ^ data_in[307] ^ data_in[305] ^ data_in[303] ^ data_in[301] ^ data_in[299] ^ data_in[297] ^ data_in[295] ^ data_in[293] ^ data_in[291] ^ data_in[289] ^ data_in[287] ^ data_in[285] ^ data_in[283] ^ data_in[281] ^ data_in[279] ^ data_in[277] ^ data_in[275] ^ data_in[273] ^ data_in[271] ^ data_in[269] ^ data_in[267] ^ data_in[265] ^ data_in[263] ^ data_in[261] ^ data_in[259] ^ data_in[257] ^ data_in[255] ^ data_in[254] ^ data_in[252] ^ data_in[250] ^ data_in[248] ^ data_in[246] ^ data_in[244] ^ data_in[242] ^ data_in[240] ^ data_in[238] ^ data_in[236] ^ data_in[234] ^ data_in[232] ^ data_in[230] ^ data_in[228] ^ data_in[226] ^ data_in[224] ^ data_in[222] ^ data_in[220] ^ data_in[218] ^ data_in[216] ^ data_in[214] ^ data_in[212] ^ data_in[210] ^ data_in[208] ^ data_in[206] ^ data_in[204] ^ data_in[202] ^ data_in[200] ^ data_in[198] ^ data_in[196] ^ data_in[194] ^ data_in[192] ^ data_in[190] ^ data_in[188] ^ data_in[186] ^ data_in[184] ^ data_in[182] ^ data_in[180] ^ data_in[178] ^ data_in[176] ^ data_in[174] ^ data_in[172] ^ data_in[170] ^ data_in[168] ^ data_in[166] ^ data_in[164] ^ data_in[162] ^ data_in[160] ^ data_in[158] ^ data_in[156] ^ data_in[154] ^ data_in[152] ^ data_in[150] ^ data_in[148] ^ data_in[146] ^ data_in[144] ^ data_in[142] ^ data_in[140] ^ data_in[138] ^ data_in[136] ^ data_in[134] ^ data_in[132] ^ data_in[130] ^ data_in[128] ^ data_in[126] ^ data_in[124] ^ data_in[122] ^ data_in[120] ^ data_in[118] ^ data_in[116] ^ data_in[114] ^ data_in[112] ^ data_in[110] ^ data_in[108] ^ data_in[106] ^ data_in[104] ^ data_in[102] ^ data_in[100] ^ data_in[98] ^ data_in[96] ^ data_in[94] ^ data_in[92] ^ data_in[90] ^ data_in[88] ^ data_in[86] ^ data_in[84] ^ data_in[82] ^ data_in[80] ^ data_in[78] ^ data_in[76] ^ data_in[74] ^ data_in[72] ^ data_in[70] ^ data_in[68] ^ data_in[66] ^ data_in[64] ^ data_in[62] ^ data_in[60] ^ data_in[58] ^ data_in[56] ^ data_in[54] ^ data_in[52] ^ data_in[50] ^ data_in[48] ^ data_in[46] ^ data_in[44] ^ data_in[42] ^ data_in[40] ^ data_in[38] ^ data_in[36] ^ data_in[34] ^ data_in[32] ^ data_in[30] ^ data_in[28] ^ data_in[26] ^ data_in[24] ^ data_in[22] ^ data_in[20] ^ data_in[18] ^ data_in[16] ^ data_in[14] ^ data_in[12] ^ data_in[10] ^ data_in[8] ^ data_in[6] ^ data_in[4] ^ data_in[2] ^ data_in[0] ;
    checker_in[1] = data_in[501] ^ data_in[499] ^ data_in[498] ^ data_in[496] ^ data_in[495] ^ data_in[492] ^ data_in[491] ^ data_in[489] ^ data_in[488] ^ data_in[485] ^ data_in[484] ^ data_in[481] ^ data_in[480] ^ data_in[477] ^ data_in[476] ^ data_in[474] ^ data_in[473] ^ data_in[470] ^ data_in[469] ^ data_in[466] ^ data_in[465] ^ data_in[462] ^ data_in[461] ^ data_in[458] ^ data_in[457] ^ data_in[454] ^ data_in[453] ^ data_in[450] ^ data_in[449] ^ data_in[446] ^ data_in[445] ^ data_in[443] ^ data_in[442] ^ data_in[439] ^ data_in[438] ^ data_in[435] ^ data_in[434] ^ data_in[431] ^ data_in[430] ^ data_in[427] ^ data_in[426] ^ data_in[423] ^ data_in[422] ^ data_in[419] ^ data_in[418] ^ data_in[415] ^ data_in[414] ^ data_in[411] ^ data_in[410] ^ data_in[407] ^ data_in[406] ^ data_in[403] ^ data_in[402] ^ data_in[399] ^ data_in[398] ^ data_in[395] ^ data_in[394] ^ data_in[391] ^ data_in[390] ^ data_in[387] ^ data_in[386] ^ data_in[383] ^ data_in[382] ^ data_in[380] ^ data_in[379] ^ data_in[376] ^ data_in[375] ^ data_in[372] ^ data_in[371] ^ data_in[368] ^ data_in[367] ^ data_in[364] ^ data_in[363] ^ data_in[360] ^ data_in[359] ^ data_in[356] ^ data_in[355] ^ data_in[352] ^ data_in[351] ^ data_in[348] ^ data_in[347] ^ data_in[344] ^ data_in[343] ^ data_in[340] ^ data_in[339] ^ data_in[336] ^ data_in[335] ^ data_in[332] ^ data_in[331] ^ data_in[328] ^ data_in[327] ^ data_in[324] ^ data_in[323] ^ data_in[320] ^ data_in[319] ^ data_in[316] ^ data_in[315] ^ data_in[312] ^ data_in[311] ^ data_in[308] ^ data_in[307] ^ data_in[304] ^ data_in[303] ^ data_in[300] ^ data_in[299] ^ data_in[296] ^ data_in[295] ^ data_in[292] ^ data_in[291] ^ data_in[288] ^ data_in[287] ^ data_in[284] ^ data_in[283] ^ data_in[280] ^ data_in[279] ^ data_in[276] ^ data_in[275] ^ data_in[272] ^ data_in[271] ^ data_in[268] ^ data_in[267] ^ data_in[264] ^ data_in[263] ^ data_in[260] ^ data_in[259] ^ data_in[256] ^ data_in[255] ^ data_in[253] ^ data_in[252] ^ data_in[249] ^ data_in[248] ^ data_in[245] ^ data_in[244] ^ data_in[241] ^ data_in[240] ^ data_in[237] ^ data_in[236] ^ data_in[233] ^ data_in[232] ^ data_in[229] ^ data_in[228] ^ data_in[225] ^ data_in[224] ^ data_in[221] ^ data_in[220] ^ data_in[217] ^ data_in[216] ^ data_in[213] ^ data_in[212] ^ data_in[209] ^ data_in[208] ^ data_in[205] ^ data_in[204] ^ data_in[201] ^ data_in[200] ^ data_in[197] ^ data_in[196] ^ data_in[193] ^ data_in[192] ^ data_in[189] ^ data_in[188] ^ data_in[185] ^ data_in[184] ^ data_in[181] ^ data_in[180] ^ data_in[177] ^ data_in[176] ^ data_in[173] ^ data_in[172] ^ data_in[169] ^ data_in[168] ^ data_in[165] ^ data_in[164] ^ data_in[161] ^ data_in[160] ^ data_in[157] ^ data_in[156] ^ data_in[153] ^ data_in[152] ^ data_in[149] ^ data_in[148] ^ data_in[145] ^ data_in[144] ^ data_in[141] ^ data_in[140] ^ data_in[137] ^ data_in[136] ^ data_in[133] ^ data_in[132] ^ data_in[129] ^ data_in[128] ^ data_in[125] ^ data_in[124] ^ data_in[121] ^ data_in[120] ^ data_in[117] ^ data_in[116] ^ data_in[113] ^ data_in[112] ^ data_in[109] ^ data_in[108] ^ data_in[105] ^ data_in[104] ^ data_in[101] ^ data_in[100] ^ data_in[97] ^ data_in[96] ^ data_in[93] ^ data_in[92] ^ data_in[89] ^ data_in[88] ^ data_in[85] ^ data_in[84] ^ data_in[81] ^ data_in[80] ^ data_in[77] ^ data_in[76] ^ data_in[73] ^ data_in[72] ^ data_in[69] ^ data_in[68] ^ data_in[65] ^ data_in[64] ^ data_in[61] ^ data_in[60] ^ data_in[57] ^ data_in[56] ^ data_in[53] ^ data_in[52] ^ data_in[49] ^ data_in[48] ^ data_in[45] ^ data_in[44] ^ data_in[41] ^ data_in[40] ^ data_in[37] ^ data_in[36] ^ data_in[33] ^ data_in[32] ^ data_in[29] ^ data_in[28] ^ data_in[25] ^ data_in[24] ^ data_in[21] ^ data_in[20] ^ data_in[17] ^ data_in[16] ^ data_in[13] ^ data_in[12] ^ data_in[9] ^ data_in[8] ^ data_in[5] ^ data_in[4] ^ data_in[1] ^ data_in[0] ;
    checker_in[2] = data_in[500] ^ data_in[499] ^ data_in[498] ^ data_in[494] ^ data_in[493] ^ data_in[492] ^ data_in[491] ^ data_in[487] ^ data_in[486] ^ data_in[485] ^ data_in[484] ^ data_in[479] ^ data_in[478] ^ data_in[477] ^ data_in[476] ^ data_in[472] ^ data_in[471] ^ data_in[470] ^ data_in[469] ^ data_in[464] ^ data_in[463] ^ data_in[462] ^ data_in[461] ^ data_in[456] ^ data_in[455] ^ data_in[454] ^ data_in[453] ^ data_in[448] ^ data_in[447] ^ data_in[446] ^ data_in[445] ^ data_in[441] ^ data_in[440] ^ data_in[439] ^ data_in[438] ^ data_in[433] ^ data_in[432] ^ data_in[431] ^ data_in[430] ^ data_in[425] ^ data_in[424] ^ data_in[423] ^ data_in[422] ^ data_in[417] ^ data_in[416] ^ data_in[415] ^ data_in[414] ^ data_in[409] ^ data_in[408] ^ data_in[407] ^ data_in[406] ^ data_in[401] ^ data_in[400] ^ data_in[399] ^ data_in[398] ^ data_in[393] ^ data_in[392] ^ data_in[391] ^ data_in[390] ^ data_in[385] ^ data_in[384] ^ data_in[383] ^ data_in[382] ^ data_in[378] ^ data_in[377] ^ data_in[376] ^ data_in[375] ^ data_in[370] ^ data_in[369] ^ data_in[368] ^ data_in[367] ^ data_in[362] ^ data_in[361] ^ data_in[360] ^ data_in[359] ^ data_in[354] ^ data_in[353] ^ data_in[352] ^ data_in[351] ^ data_in[346] ^ data_in[345] ^ data_in[344] ^ data_in[343] ^ data_in[338] ^ data_in[337] ^ data_in[336] ^ data_in[335] ^ data_in[330] ^ data_in[329] ^ data_in[328] ^ data_in[327] ^ data_in[322] ^ data_in[321] ^ data_in[320] ^ data_in[319] ^ data_in[314] ^ data_in[313] ^ data_in[312] ^ data_in[311] ^ data_in[306] ^ data_in[305] ^ data_in[304] ^ data_in[303] ^ data_in[298] ^ data_in[297] ^ data_in[296] ^ data_in[295] ^ data_in[290] ^ data_in[289] ^ data_in[288] ^ data_in[287] ^ data_in[282] ^ data_in[281] ^ data_in[280] ^ data_in[279] ^ data_in[274] ^ data_in[273] ^ data_in[272] ^ data_in[271] ^ data_in[266] ^ data_in[265] ^ data_in[264] ^ data_in[263] ^ data_in[258] ^ data_in[257] ^ data_in[256] ^ data_in[255] ^ data_in[251] ^ data_in[250] ^ data_in[249] ^ data_in[248] ^ data_in[243] ^ data_in[242] ^ data_in[241] ^ data_in[240] ^ data_in[235] ^ data_in[234] ^ data_in[233] ^ data_in[232] ^ data_in[227] ^ data_in[226] ^ data_in[225] ^ data_in[224] ^ data_in[219] ^ data_in[218] ^ data_in[217] ^ data_in[216] ^ data_in[211] ^ data_in[210] ^ data_in[209] ^ data_in[208] ^ data_in[203] ^ data_in[202] ^ data_in[201] ^ data_in[200] ^ data_in[195] ^ data_in[194] ^ data_in[193] ^ data_in[192] ^ data_in[187] ^ data_in[186] ^ data_in[185] ^ data_in[184] ^ data_in[179] ^ data_in[178] ^ data_in[177] ^ data_in[176] ^ data_in[171] ^ data_in[170] ^ data_in[169] ^ data_in[168] ^ data_in[163] ^ data_in[162] ^ data_in[161] ^ data_in[160] ^ data_in[155] ^ data_in[154] ^ data_in[153] ^ data_in[152] ^ data_in[147] ^ data_in[146] ^ data_in[145] ^ data_in[144] ^ data_in[139] ^ data_in[138] ^ data_in[137] ^ data_in[136] ^ data_in[131] ^ data_in[130] ^ data_in[129] ^ data_in[128] ^ data_in[123] ^ data_in[122] ^ data_in[121] ^ data_in[120] ^ data_in[115] ^ data_in[114] ^ data_in[113] ^ data_in[112] ^ data_in[107] ^ data_in[106] ^ data_in[105] ^ data_in[104] ^ data_in[99] ^ data_in[98] ^ data_in[97] ^ data_in[96] ^ data_in[91] ^ data_in[90] ^ data_in[89] ^ data_in[88] ^ data_in[83] ^ data_in[82] ^ data_in[81] ^ data_in[80] ^ data_in[75] ^ data_in[74] ^ data_in[73] ^ data_in[72] ^ data_in[67] ^ data_in[66] ^ data_in[65] ^ data_in[64] ^ data_in[59] ^ data_in[58] ^ data_in[57] ^ data_in[56] ^ data_in[51] ^ data_in[50] ^ data_in[49] ^ data_in[48] ^ data_in[43] ^ data_in[42] ^ data_in[41] ^ data_in[40] ^ data_in[35] ^ data_in[34] ^ data_in[33] ^ data_in[32] ^ data_in[27] ^ data_in[26] ^ data_in[25] ^ data_in[24] ^ data_in[19] ^ data_in[18] ^ data_in[17] ^ data_in[16] ^ data_in[11] ^ data_in[10] ^ data_in[9] ^ data_in[8] ^ data_in[3] ^ data_in[2] ^ data_in[1] ^ data_in[0] ;
    checker_in[3] = data_in[497] ^ data_in[496] ^ data_in[495] ^ data_in[494] ^ data_in[493] ^ data_in[492] ^ data_in[491] ^ data_in[483] ^ data_in[482] ^ data_in[481] ^ data_in[480] ^ data_in[479] ^ data_in[478] ^ data_in[477] ^ data_in[476] ^ data_in[468] ^ data_in[467] ^ data_in[466] ^ data_in[465] ^ data_in[464] ^ data_in[463] ^ data_in[462] ^ data_in[461] ^ data_in[452] ^ data_in[451] ^ data_in[450] ^ data_in[449] ^ data_in[448] ^ data_in[447] ^ data_in[446] ^ data_in[445] ^ data_in[437] ^ data_in[436] ^ data_in[435] ^ data_in[434] ^ data_in[433] ^ data_in[432] ^ data_in[431] ^ data_in[430] ^ data_in[421] ^ data_in[420] ^ data_in[419] ^ data_in[418] ^ data_in[417] ^ data_in[416] ^ data_in[415] ^ data_in[414] ^ data_in[405] ^ data_in[404] ^ data_in[403] ^ data_in[402] ^ data_in[401] ^ data_in[400] ^ data_in[399] ^ data_in[398] ^ data_in[389] ^ data_in[388] ^ data_in[387] ^ data_in[386] ^ data_in[385] ^ data_in[384] ^ data_in[383] ^ data_in[382] ^ data_in[374] ^ data_in[373] ^ data_in[372] ^ data_in[371] ^ data_in[370] ^ data_in[369] ^ data_in[368] ^ data_in[367] ^ data_in[358] ^ data_in[357] ^ data_in[356] ^ data_in[355] ^ data_in[354] ^ data_in[353] ^ data_in[352] ^ data_in[351] ^ data_in[342] ^ data_in[341] ^ data_in[340] ^ data_in[339] ^ data_in[338] ^ data_in[337] ^ data_in[336] ^ data_in[335] ^ data_in[326] ^ data_in[325] ^ data_in[324] ^ data_in[323] ^ data_in[322] ^ data_in[321] ^ data_in[320] ^ data_in[319] ^ data_in[310] ^ data_in[309] ^ data_in[308] ^ data_in[307] ^ data_in[306] ^ data_in[305] ^ data_in[304] ^ data_in[303] ^ data_in[294] ^ data_in[293] ^ data_in[292] ^ data_in[291] ^ data_in[290] ^ data_in[289] ^ data_in[288] ^ data_in[287] ^ data_in[278] ^ data_in[277] ^ data_in[276] ^ data_in[275] ^ data_in[274] ^ data_in[273] ^ data_in[272] ^ data_in[271] ^ data_in[262] ^ data_in[261] ^ data_in[260] ^ data_in[259] ^ data_in[258] ^ data_in[257] ^ data_in[256] ^ data_in[255] ^ data_in[247] ^ data_in[246] ^ data_in[245] ^ data_in[244] ^ data_in[243] ^ data_in[242] ^ data_in[241] ^ data_in[240] ^ data_in[231] ^ data_in[230] ^ data_in[229] ^ data_in[228] ^ data_in[227] ^ data_in[226] ^ data_in[225] ^ data_in[224] ^ data_in[215] ^ data_in[214] ^ data_in[213] ^ data_in[212] ^ data_in[211] ^ data_in[210] ^ data_in[209] ^ data_in[208] ^ data_in[199] ^ data_in[198] ^ data_in[197] ^ data_in[196] ^ data_in[195] ^ data_in[194] ^ data_in[193] ^ data_in[192] ^ data_in[183] ^ data_in[182] ^ data_in[181] ^ data_in[180] ^ data_in[179] ^ data_in[178] ^ data_in[177] ^ data_in[176] ^ data_in[167] ^ data_in[166] ^ data_in[165] ^ data_in[164] ^ data_in[163] ^ data_in[162] ^ data_in[161] ^ data_in[160] ^ data_in[151] ^ data_in[150] ^ data_in[149] ^ data_in[148] ^ data_in[147] ^ data_in[146] ^ data_in[145] ^ data_in[144] ^ data_in[135] ^ data_in[134] ^ data_in[133] ^ data_in[132] ^ data_in[131] ^ data_in[130] ^ data_in[129] ^ data_in[128] ^ data_in[119] ^ data_in[118] ^ data_in[117] ^ data_in[116] ^ data_in[115] ^ data_in[114] ^ data_in[113] ^ data_in[112] ^ data_in[103] ^ data_in[102] ^ data_in[101] ^ data_in[100] ^ data_in[99] ^ data_in[98] ^ data_in[97] ^ data_in[96] ^ data_in[87] ^ data_in[86] ^ data_in[85] ^ data_in[84] ^ data_in[83] ^ data_in[82] ^ data_in[81] ^ data_in[80] ^ data_in[71] ^ data_in[70] ^ data_in[69] ^ data_in[68] ^ data_in[67] ^ data_in[66] ^ data_in[65] ^ data_in[64] ^ data_in[55] ^ data_in[54] ^ data_in[53] ^ data_in[52] ^ data_in[51] ^ data_in[50] ^ data_in[49] ^ data_in[48] ^ data_in[39] ^ data_in[38] ^ data_in[37] ^ data_in[36] ^ data_in[35] ^ data_in[34] ^ data_in[33] ^ data_in[32] ^ data_in[23] ^ data_in[22] ^ data_in[21] ^ data_in[20] ^ data_in[19] ^ data_in[18] ^ data_in[17] ^ data_in[16] ^ data_in[7] ^ data_in[6] ^ data_in[5] ^ data_in[4] ^ data_in[3] ^ data_in[2] ^ data_in[1] ^ data_in[0] ;
    checker_in[4] = data_in[490] ^ data_in[489] ^ data_in[488] ^ data_in[487] ^ data_in[486] ^ data_in[485] ^ data_in[484] ^ data_in[483] ^ data_in[482] ^ data_in[481] ^ data_in[480] ^ data_in[479] ^ data_in[478] ^ data_in[477] ^ data_in[476] ^ data_in[460] ^ data_in[459] ^ data_in[458] ^ data_in[457] ^ data_in[456] ^ data_in[455] ^ data_in[454] ^ data_in[453] ^ data_in[452] ^ data_in[451] ^ data_in[450] ^ data_in[449] ^ data_in[448] ^ data_in[447] ^ data_in[446] ^ data_in[445] ^ data_in[429] ^ data_in[428] ^ data_in[427] ^ data_in[426] ^ data_in[425] ^ data_in[424] ^ data_in[423] ^ data_in[422] ^ data_in[421] ^ data_in[420] ^ data_in[419] ^ data_in[418] ^ data_in[417] ^ data_in[416] ^ data_in[415] ^ data_in[414] ^ data_in[397] ^ data_in[396] ^ data_in[395] ^ data_in[394] ^ data_in[393] ^ data_in[392] ^ data_in[391] ^ data_in[390] ^ data_in[389] ^ data_in[388] ^ data_in[387] ^ data_in[386] ^ data_in[385] ^ data_in[384] ^ data_in[383] ^ data_in[382] ^ data_in[366] ^ data_in[365] ^ data_in[364] ^ data_in[363] ^ data_in[362] ^ data_in[361] ^ data_in[360] ^ data_in[359] ^ data_in[358] ^ data_in[357] ^ data_in[356] ^ data_in[355] ^ data_in[354] ^ data_in[353] ^ data_in[352] ^ data_in[351] ^ data_in[334] ^ data_in[333] ^ data_in[332] ^ data_in[331] ^ data_in[330] ^ data_in[329] ^ data_in[328] ^ data_in[327] ^ data_in[326] ^ data_in[325] ^ data_in[324] ^ data_in[323] ^ data_in[322] ^ data_in[321] ^ data_in[320] ^ data_in[319] ^ data_in[302] ^ data_in[301] ^ data_in[300] ^ data_in[299] ^ data_in[298] ^ data_in[297] ^ data_in[296] ^ data_in[295] ^ data_in[294] ^ data_in[293] ^ data_in[292] ^ data_in[291] ^ data_in[290] ^ data_in[289] ^ data_in[288] ^ data_in[287] ^ data_in[270] ^ data_in[269] ^ data_in[268] ^ data_in[267] ^ data_in[266] ^ data_in[265] ^ data_in[264] ^ data_in[263] ^ data_in[262] ^ data_in[261] ^ data_in[260] ^ data_in[259] ^ data_in[258] ^ data_in[257] ^ data_in[256] ^ data_in[255] ^ data_in[239] ^ data_in[238] ^ data_in[237] ^ data_in[236] ^ data_in[235] ^ data_in[234] ^ data_in[233] ^ data_in[232] ^ data_in[231] ^ data_in[230] ^ data_in[229] ^ data_in[228] ^ data_in[227] ^ data_in[226] ^ data_in[225] ^ data_in[224] ^ data_in[207] ^ data_in[206] ^ data_in[205] ^ data_in[204] ^ data_in[203] ^ data_in[202] ^ data_in[201] ^ data_in[200] ^ data_in[199] ^ data_in[198] ^ data_in[197] ^ data_in[196] ^ data_in[195] ^ data_in[194] ^ data_in[193] ^ data_in[192] ^ data_in[175] ^ data_in[174] ^ data_in[173] ^ data_in[172] ^ data_in[171] ^ data_in[170] ^ data_in[169] ^ data_in[168] ^ data_in[167] ^ data_in[166] ^ data_in[165] ^ data_in[164] ^ data_in[163] ^ data_in[162] ^ data_in[161] ^ data_in[160] ^ data_in[143] ^ data_in[142] ^ data_in[141] ^ data_in[140] ^ data_in[139] ^ data_in[138] ^ data_in[137] ^ data_in[136] ^ data_in[135] ^ data_in[134] ^ data_in[133] ^ data_in[132] ^ data_in[131] ^ data_in[130] ^ data_in[129] ^ data_in[128] ^ data_in[111] ^ data_in[110] ^ data_in[109] ^ data_in[108] ^ data_in[107] ^ data_in[106] ^ data_in[105] ^ data_in[104] ^ data_in[103] ^ data_in[102] ^ data_in[101] ^ data_in[100] ^ data_in[99] ^ data_in[98] ^ data_in[97] ^ data_in[96] ^ data_in[79] ^ data_in[78] ^ data_in[77] ^ data_in[76] ^ data_in[75] ^ data_in[74] ^ data_in[73] ^ data_in[72] ^ data_in[71] ^ data_in[70] ^ data_in[69] ^ data_in[68] ^ data_in[67] ^ data_in[66] ^ data_in[65] ^ data_in[64] ^ data_in[47] ^ data_in[46] ^ data_in[45] ^ data_in[44] ^ data_in[43] ^ data_in[42] ^ data_in[41] ^ data_in[40] ^ data_in[39] ^ data_in[38] ^ data_in[37] ^ data_in[36] ^ data_in[35] ^ data_in[34] ^ data_in[33] ^ data_in[32] ^ data_in[15] ^ data_in[14] ^ data_in[13] ^ data_in[12] ^ data_in[11] ^ data_in[10] ^ data_in[9] ^ data_in[8] ^ data_in[7] ^ data_in[6] ^ data_in[5] ^ data_in[4] ^ data_in[3] ^ data_in[2] ^ data_in[1] ^ data_in[0] ;
    checker_in[5] = data_in[475] ^ data_in[474] ^ data_in[473] ^ data_in[472] ^ data_in[471] ^ data_in[470] ^ data_in[469] ^ data_in[468] ^ data_in[467] ^ data_in[466] ^ data_in[465] ^ data_in[464] ^ data_in[463] ^ data_in[462] ^ data_in[461] ^ data_in[460] ^ data_in[459] ^ data_in[458] ^ data_in[457] ^ data_in[456] ^ data_in[455] ^ data_in[454] ^ data_in[453] ^ data_in[452] ^ data_in[451] ^ data_in[450] ^ data_in[449] ^ data_in[448] ^ data_in[447] ^ data_in[446] ^ data_in[445] ^ data_in[413] ^ data_in[412] ^ data_in[411] ^ data_in[410] ^ data_in[409] ^ data_in[408] ^ data_in[407] ^ data_in[406] ^ data_in[405] ^ data_in[404] ^ data_in[403] ^ data_in[402] ^ data_in[401] ^ data_in[400] ^ data_in[399] ^ data_in[398] ^ data_in[397] ^ data_in[396] ^ data_in[395] ^ data_in[394] ^ data_in[393] ^ data_in[392] ^ data_in[391] ^ data_in[390] ^ data_in[389] ^ data_in[388] ^ data_in[387] ^ data_in[386] ^ data_in[385] ^ data_in[384] ^ data_in[383] ^ data_in[382] ^ data_in[350] ^ data_in[349] ^ data_in[348] ^ data_in[347] ^ data_in[346] ^ data_in[345] ^ data_in[344] ^ data_in[343] ^ data_in[342] ^ data_in[341] ^ data_in[340] ^ data_in[339] ^ data_in[338] ^ data_in[337] ^ data_in[336] ^ data_in[335] ^ data_in[334] ^ data_in[333] ^ data_in[332] ^ data_in[331] ^ data_in[330] ^ data_in[329] ^ data_in[328] ^ data_in[327] ^ data_in[326] ^ data_in[325] ^ data_in[324] ^ data_in[323] ^ data_in[322] ^ data_in[321] ^ data_in[320] ^ data_in[319] ^ data_in[286] ^ data_in[285] ^ data_in[284] ^ data_in[283] ^ data_in[282] ^ data_in[281] ^ data_in[280] ^ data_in[279] ^ data_in[278] ^ data_in[277] ^ data_in[276] ^ data_in[275] ^ data_in[274] ^ data_in[273] ^ data_in[272] ^ data_in[271] ^ data_in[270] ^ data_in[269] ^ data_in[268] ^ data_in[267] ^ data_in[266] ^ data_in[265] ^ data_in[264] ^ data_in[263] ^ data_in[262] ^ data_in[261] ^ data_in[260] ^ data_in[259] ^ data_in[258] ^ data_in[257] ^ data_in[256] ^ data_in[255] ^ data_in[223] ^ data_in[222] ^ data_in[221] ^ data_in[220] ^ data_in[219] ^ data_in[218] ^ data_in[217] ^ data_in[216] ^ data_in[215] ^ data_in[214] ^ data_in[213] ^ data_in[212] ^ data_in[211] ^ data_in[210] ^ data_in[209] ^ data_in[208] ^ data_in[207] ^ data_in[206] ^ data_in[205] ^ data_in[204] ^ data_in[203] ^ data_in[202] ^ data_in[201] ^ data_in[200] ^ data_in[199] ^ data_in[198] ^ data_in[197] ^ data_in[196] ^ data_in[195] ^ data_in[194] ^ data_in[193] ^ data_in[192] ^ data_in[159] ^ data_in[158] ^ data_in[157] ^ data_in[156] ^ data_in[155] ^ data_in[154] ^ data_in[153] ^ data_in[152] ^ data_in[151] ^ data_in[150] ^ data_in[149] ^ data_in[148] ^ data_in[147] ^ data_in[146] ^ data_in[145] ^ data_in[144] ^ data_in[143] ^ data_in[142] ^ data_in[141] ^ data_in[140] ^ data_in[139] ^ data_in[138] ^ data_in[137] ^ data_in[136] ^ data_in[135] ^ data_in[134] ^ data_in[133] ^ data_in[132] ^ data_in[131] ^ data_in[130] ^ data_in[129] ^ data_in[128] ^ data_in[95] ^ data_in[94] ^ data_in[93] ^ data_in[92] ^ data_in[91] ^ data_in[90] ^ data_in[89] ^ data_in[88] ^ data_in[87] ^ data_in[86] ^ data_in[85] ^ data_in[84] ^ data_in[83] ^ data_in[82] ^ data_in[81] ^ data_in[80] ^ data_in[79] ^ data_in[78] ^ data_in[77] ^ data_in[76] ^ data_in[75] ^ data_in[74] ^ data_in[73] ^ data_in[72] ^ data_in[71] ^ data_in[70] ^ data_in[69] ^ data_in[68] ^ data_in[67] ^ data_in[66] ^ data_in[65] ^ data_in[64] ^ data_in[31] ^ data_in[30] ^ data_in[29] ^ data_in[28] ^ data_in[27] ^ data_in[26] ^ data_in[25] ^ data_in[24] ^ data_in[23] ^ data_in[22] ^ data_in[21] ^ data_in[20] ^ data_in[19] ^ data_in[18] ^ data_in[17] ^ data_in[16] ^ data_in[15] ^ data_in[14] ^ data_in[13] ^ data_in[12] ^ data_in[11] ^ data_in[10] ^ data_in[9] ^ data_in[8] ^ data_in[7] ^ data_in[6] ^ data_in[5] ^ data_in[4] ^ data_in[3] ^ data_in[2] ^ data_in[1] ^ data_in[0] ;
    checker_in[6] = data_in[444] ^ data_in[443] ^ data_in[442] ^ data_in[441] ^ data_in[440] ^ data_in[439] ^ data_in[438] ^ data_in[437] ^ data_in[436] ^ data_in[435] ^ data_in[434] ^ data_in[433] ^ data_in[432] ^ data_in[431] ^ data_in[430] ^ data_in[429] ^ data_in[428] ^ data_in[427] ^ data_in[426] ^ data_in[425] ^ data_in[424] ^ data_in[423] ^ data_in[422] ^ data_in[421] ^ data_in[420] ^ data_in[419] ^ data_in[418] ^ data_in[417] ^ data_in[416] ^ data_in[415] ^ data_in[414] ^ data_in[413] ^ data_in[412] ^ data_in[411] ^ data_in[410] ^ data_in[409] ^ data_in[408] ^ data_in[407] ^ data_in[406] ^ data_in[405] ^ data_in[404] ^ data_in[403] ^ data_in[402] ^ data_in[401] ^ data_in[400] ^ data_in[399] ^ data_in[398] ^ data_in[397] ^ data_in[396] ^ data_in[395] ^ data_in[394] ^ data_in[393] ^ data_in[392] ^ data_in[391] ^ data_in[390] ^ data_in[389] ^ data_in[388] ^ data_in[387] ^ data_in[386] ^ data_in[385] ^ data_in[384] ^ data_in[383] ^ data_in[382] ^ data_in[318] ^ data_in[317] ^ data_in[316] ^ data_in[315] ^ data_in[314] ^ data_in[313] ^ data_in[312] ^ data_in[311] ^ data_in[310] ^ data_in[309] ^ data_in[308] ^ data_in[307] ^ data_in[306] ^ data_in[305] ^ data_in[304] ^ data_in[303] ^ data_in[302] ^ data_in[301] ^ data_in[300] ^ data_in[299] ^ data_in[298] ^ data_in[297] ^ data_in[296] ^ data_in[295] ^ data_in[294] ^ data_in[293] ^ data_in[292] ^ data_in[291] ^ data_in[290] ^ data_in[289] ^ data_in[288] ^ data_in[287] ^ data_in[286] ^ data_in[285] ^ data_in[284] ^ data_in[283] ^ data_in[282] ^ data_in[281] ^ data_in[280] ^ data_in[279] ^ data_in[278] ^ data_in[277] ^ data_in[276] ^ data_in[275] ^ data_in[274] ^ data_in[273] ^ data_in[272] ^ data_in[271] ^ data_in[270] ^ data_in[269] ^ data_in[268] ^ data_in[267] ^ data_in[266] ^ data_in[265] ^ data_in[264] ^ data_in[263] ^ data_in[262] ^ data_in[261] ^ data_in[260] ^ data_in[259] ^ data_in[258] ^ data_in[257] ^ data_in[256] ^ data_in[255] ^ data_in[191] ^ data_in[190] ^ data_in[189] ^ data_in[188] ^ data_in[187] ^ data_in[186] ^ data_in[185] ^ data_in[184] ^ data_in[183] ^ data_in[182] ^ data_in[181] ^ data_in[180] ^ data_in[179] ^ data_in[178] ^ data_in[177] ^ data_in[176] ^ data_in[175] ^ data_in[174] ^ data_in[173] ^ data_in[172] ^ data_in[171] ^ data_in[170] ^ data_in[169] ^ data_in[168] ^ data_in[167] ^ data_in[166] ^ data_in[165] ^ data_in[164] ^ data_in[163] ^ data_in[162] ^ data_in[161] ^ data_in[160] ^ data_in[159] ^ data_in[158] ^ data_in[157] ^ data_in[156] ^ data_in[155] ^ data_in[154] ^ data_in[153] ^ data_in[152] ^ data_in[151] ^ data_in[150] ^ data_in[149] ^ data_in[148] ^ data_in[147] ^ data_in[146] ^ data_in[145] ^ data_in[144] ^ data_in[143] ^ data_in[142] ^ data_in[141] ^ data_in[140] ^ data_in[139] ^ data_in[138] ^ data_in[137] ^ data_in[136] ^ data_in[135] ^ data_in[134] ^ data_in[133] ^ data_in[132] ^ data_in[131] ^ data_in[130] ^ data_in[129] ^ data_in[128] ^ data_in[63] ^ data_in[62] ^ data_in[61] ^ data_in[60] ^ data_in[59] ^ data_in[58] ^ data_in[57] ^ data_in[56] ^ data_in[55] ^ data_in[54] ^ data_in[53] ^ data_in[52] ^ data_in[51] ^ data_in[50] ^ data_in[49] ^ data_in[48] ^ data_in[47] ^ data_in[46] ^ data_in[45] ^ data_in[44] ^ data_in[43] ^ data_in[42] ^ data_in[41] ^ data_in[40] ^ data_in[39] ^ data_in[38] ^ data_in[37] ^ data_in[36] ^ data_in[35] ^ data_in[34] ^ data_in[33] ^ data_in[32] ^ data_in[31] ^ data_in[30] ^ data_in[29] ^ data_in[28] ^ data_in[27] ^ data_in[26] ^ data_in[25] ^ data_in[24] ^ data_in[23] ^ data_in[22] ^ data_in[21] ^ data_in[20] ^ data_in[19] ^ data_in[18] ^ data_in[17] ^ data_in[16] ^ data_in[15] ^ data_in[14] ^ data_in[13] ^ data_in[12] ^ data_in[11] ^ data_in[10] ^ data_in[9] ^ data_in[8] ^ data_in[7] ^ data_in[6] ^ data_in[5] ^ data_in[4] ^ data_in[3] ^ data_in[2] ^ data_in[1] ^ data_in[0] ;
    checker_in[7] = data_in[381] ^ data_in[380] ^ data_in[379] ^ data_in[378] ^ data_in[377] ^ data_in[376] ^ data_in[375] ^ data_in[374] ^ data_in[373] ^ data_in[372] ^ data_in[371] ^ data_in[370] ^ data_in[369] ^ data_in[368] ^ data_in[367] ^ data_in[366] ^ data_in[365] ^ data_in[364] ^ data_in[363] ^ data_in[362] ^ data_in[361] ^ data_in[360] ^ data_in[359] ^ data_in[358] ^ data_in[357] ^ data_in[356] ^ data_in[355] ^ data_in[354] ^ data_in[353] ^ data_in[352] ^ data_in[351] ^ data_in[350] ^ data_in[349] ^ data_in[348] ^ data_in[347] ^ data_in[346] ^ data_in[345] ^ data_in[344] ^ data_in[343] ^ data_in[342] ^ data_in[341] ^ data_in[340] ^ data_in[339] ^ data_in[338] ^ data_in[337] ^ data_in[336] ^ data_in[335] ^ data_in[334] ^ data_in[333] ^ data_in[332] ^ data_in[331] ^ data_in[330] ^ data_in[329] ^ data_in[328] ^ data_in[327] ^ data_in[326] ^ data_in[325] ^ data_in[324] ^ data_in[323] ^ data_in[322] ^ data_in[321] ^ data_in[320] ^ data_in[319] ^ data_in[318] ^ data_in[317] ^ data_in[316] ^ data_in[315] ^ data_in[314] ^ data_in[313] ^ data_in[312] ^ data_in[311] ^ data_in[310] ^ data_in[309] ^ data_in[308] ^ data_in[307] ^ data_in[306] ^ data_in[305] ^ data_in[304] ^ data_in[303] ^ data_in[302] ^ data_in[301] ^ data_in[300] ^ data_in[299] ^ data_in[298] ^ data_in[297] ^ data_in[296] ^ data_in[295] ^ data_in[294] ^ data_in[293] ^ data_in[292] ^ data_in[291] ^ data_in[290] ^ data_in[289] ^ data_in[288] ^ data_in[287] ^ data_in[286] ^ data_in[285] ^ data_in[284] ^ data_in[283] ^ data_in[282] ^ data_in[281] ^ data_in[280] ^ data_in[279] ^ data_in[278] ^ data_in[277] ^ data_in[276] ^ data_in[275] ^ data_in[274] ^ data_in[273] ^ data_in[272] ^ data_in[271] ^ data_in[270] ^ data_in[269] ^ data_in[268] ^ data_in[267] ^ data_in[266] ^ data_in[265] ^ data_in[264] ^ data_in[263] ^ data_in[262] ^ data_in[261] ^ data_in[260] ^ data_in[259] ^ data_in[258] ^ data_in[257] ^ data_in[256] ^ data_in[255] ^ data_in[127] ^ data_in[126] ^ data_in[125] ^ data_in[124] ^ data_in[123] ^ data_in[122] ^ data_in[121] ^ data_in[120] ^ data_in[119] ^ data_in[118] ^ data_in[117] ^ data_in[116] ^ data_in[115] ^ data_in[114] ^ data_in[113] ^ data_in[112] ^ data_in[111] ^ data_in[110] ^ data_in[109] ^ data_in[108] ^ data_in[107] ^ data_in[106] ^ data_in[105] ^ data_in[104] ^ data_in[103] ^ data_in[102] ^ data_in[101] ^ data_in[100] ^ data_in[99] ^ data_in[98] ^ data_in[97] ^ data_in[96] ^ data_in[95] ^ data_in[94] ^ data_in[93] ^ data_in[92] ^ data_in[91] ^ data_in[90] ^ data_in[89] ^ data_in[88] ^ data_in[87] ^ data_in[86] ^ data_in[85] ^ data_in[84] ^ data_in[83] ^ data_in[82] ^ data_in[81] ^ data_in[80] ^ data_in[79] ^ data_in[78] ^ data_in[77] ^ data_in[76] ^ data_in[75] ^ data_in[74] ^ data_in[73] ^ data_in[72] ^ data_in[71] ^ data_in[70] ^ data_in[69] ^ data_in[68] ^ data_in[67] ^ data_in[66] ^ data_in[65] ^ data_in[64] ^ data_in[63] ^ data_in[62] ^ data_in[61] ^ data_in[60] ^ data_in[59] ^ data_in[58] ^ data_in[57] ^ data_in[56] ^ data_in[55] ^ data_in[54] ^ data_in[53] ^ data_in[52] ^ data_in[51] ^ data_in[50] ^ data_in[49] ^ data_in[48] ^ data_in[47] ^ data_in[46] ^ data_in[45] ^ data_in[44] ^ data_in[43] ^ data_in[42] ^ data_in[41] ^ data_in[40] ^ data_in[39] ^ data_in[38] ^ data_in[37] ^ data_in[36] ^ data_in[35] ^ data_in[34] ^ data_in[33] ^ data_in[32] ^ data_in[31] ^ data_in[30] ^ data_in[29] ^ data_in[28] ^ data_in[27] ^ data_in[26] ^ data_in[25] ^ data_in[24] ^ data_in[23] ^ data_in[22] ^ data_in[21] ^ data_in[20] ^ data_in[19] ^ data_in[18] ^ data_in[17] ^ data_in[16] ^ data_in[15] ^ data_in[14] ^ data_in[13] ^ data_in[12] ^ data_in[11] ^ data_in[10] ^ data_in[9] ^ data_in[8] ^ data_in[7] ^ data_in[6] ^ data_in[5] ^ data_in[4] ^ data_in[3] ^ data_in[2] ^ data_in[1] ^ data_in[0] ;
    checker_in[8] = data_in[254] ^ data_in[253] ^ data_in[252] ^ data_in[251] ^ data_in[250] ^ data_in[249] ^ data_in[248] ^ data_in[247] ^ data_in[246] ^ data_in[245] ^ data_in[244] ^ data_in[243] ^ data_in[242] ^ data_in[241] ^ data_in[240] ^ data_in[239] ^ data_in[238] ^ data_in[237] ^ data_in[236] ^ data_in[235] ^ data_in[234] ^ data_in[233] ^ data_in[232] ^ data_in[231] ^ data_in[230] ^ data_in[229] ^ data_in[228] ^ data_in[227] ^ data_in[226] ^ data_in[225] ^ data_in[224] ^ data_in[223] ^ data_in[222] ^ data_in[221] ^ data_in[220] ^ data_in[219] ^ data_in[218] ^ data_in[217] ^ data_in[216] ^ data_in[215] ^ data_in[214] ^ data_in[213] ^ data_in[212] ^ data_in[211] ^ data_in[210] ^ data_in[209] ^ data_in[208] ^ data_in[207] ^ data_in[206] ^ data_in[205] ^ data_in[204] ^ data_in[203] ^ data_in[202] ^ data_in[201] ^ data_in[200] ^ data_in[199] ^ data_in[198] ^ data_in[197] ^ data_in[196] ^ data_in[195] ^ data_in[194] ^ data_in[193] ^ data_in[192] ^ data_in[191] ^ data_in[190] ^ data_in[189] ^ data_in[188] ^ data_in[187] ^ data_in[186] ^ data_in[185] ^ data_in[184] ^ data_in[183] ^ data_in[182] ^ data_in[181] ^ data_in[180] ^ data_in[179] ^ data_in[178] ^ data_in[177] ^ data_in[176] ^ data_in[175] ^ data_in[174] ^ data_in[173] ^ data_in[172] ^ data_in[171] ^ data_in[170] ^ data_in[169] ^ data_in[168] ^ data_in[167] ^ data_in[166] ^ data_in[165] ^ data_in[164] ^ data_in[163] ^ data_in[162] ^ data_in[161] ^ data_in[160] ^ data_in[159] ^ data_in[158] ^ data_in[157] ^ data_in[156] ^ data_in[155] ^ data_in[154] ^ data_in[153] ^ data_in[152] ^ data_in[151] ^ data_in[150] ^ data_in[149] ^ data_in[148] ^ data_in[147] ^ data_in[146] ^ data_in[145] ^ data_in[144] ^ data_in[143] ^ data_in[142] ^ data_in[141] ^ data_in[140] ^ data_in[139] ^ data_in[138] ^ data_in[137] ^ data_in[136] ^ data_in[135] ^ data_in[134] ^ data_in[133] ^ data_in[132] ^ data_in[131] ^ data_in[130] ^ data_in[129] ^ data_in[128] ^ data_in[127] ^ data_in[126] ^ data_in[125] ^ data_in[124] ^ data_in[123] ^ data_in[122] ^ data_in[121] ^ data_in[120] ^ data_in[119] ^ data_in[118] ^ data_in[117] ^ data_in[116] ^ data_in[115] ^ data_in[114] ^ data_in[113] ^ data_in[112] ^ data_in[111] ^ data_in[110] ^ data_in[109] ^ data_in[108] ^ data_in[107] ^ data_in[106] ^ data_in[105] ^ data_in[104] ^ data_in[103] ^ data_in[102] ^ data_in[101] ^ data_in[100] ^ data_in[99] ^ data_in[98] ^ data_in[97] ^ data_in[96] ^ data_in[95] ^ data_in[94] ^ data_in[93] ^ data_in[92] ^ data_in[91] ^ data_in[90] ^ data_in[89] ^ data_in[88] ^ data_in[87] ^ data_in[86] ^ data_in[85] ^ data_in[84] ^ data_in[83] ^ data_in[82] ^ data_in[81] ^ data_in[80] ^ data_in[79] ^ data_in[78] ^ data_in[77] ^ data_in[76] ^ data_in[75] ^ data_in[74] ^ data_in[73] ^ data_in[72] ^ data_in[71] ^ data_in[70] ^ data_in[69] ^ data_in[68] ^ data_in[67] ^ data_in[66] ^ data_in[65] ^ data_in[64] ^ data_in[63] ^ data_in[62] ^ data_in[61] ^ data_in[60] ^ data_in[59] ^ data_in[58] ^ data_in[57] ^ data_in[56] ^ data_in[55] ^ data_in[54] ^ data_in[53] ^ data_in[52] ^ data_in[51] ^ data_in[50] ^ data_in[49] ^ data_in[48] ^ data_in[47] ^ data_in[46] ^ data_in[45] ^ data_in[44] ^ data_in[43] ^ data_in[42] ^ data_in[41] ^ data_in[40] ^ data_in[39] ^ data_in[38] ^ data_in[37] ^ data_in[36] ^ data_in[35] ^ data_in[34] ^ data_in[33] ^ data_in[32] ^ data_in[31] ^ data_in[30] ^ data_in[29] ^ data_in[28] ^ data_in[27] ^ data_in[26] ^ data_in[25] ^ data_in[24] ^ data_in[23] ^ data_in[22] ^ data_in[21] ^ data_in[20] ^ data_in[19] ^ data_in[18] ^ data_in[17] ^ data_in[16] ^ data_in[15] ^ data_in[14] ^ data_in[13] ^ data_in[12] ^ data_in[11] ^ data_in[10] ^ data_in[9] ^ data_in[8] ^ data_in[7] ^ data_in[6] ^ data_in[5] ^ data_in[4] ^ data_in[3] ^ data_in[2] ^ data_in[1] ^ data_in[0] ;
    parity_in = data_in[0] ^ data_in[1] ^ data_in[2] ^ data_in[3] ^ data_in[4] ^ data_in[5] ^ data_in[6] ^ data_in[7] ^ data_in[8] ^ data_in[9] ^ data_in[10] ^ data_in[11] ^ data_in[12] ^ data_in[13] ^ data_in[14] ^ data_in[15] ^ data_in[16] ^ data_in[17] ^ data_in[18] ^ data_in[19] ^ data_in[20] ^ data_in[21] ^ data_in[22] ^ data_in[23] ^ data_in[24] ^ data_in[25] ^ data_in[26] ^ data_in[27] ^ data_in[28] ^ data_in[29] ^ data_in[30] ^ data_in[31] ^ data_in[32] ^ data_in[33] ^ data_in[34] ^ data_in[35] ^ data_in[36] ^ data_in[37] ^ data_in[38] ^ data_in[39] ^ data_in[40] ^ data_in[41] ^ data_in[42] ^ data_in[43] ^ data_in[44] ^ data_in[45] ^ data_in[46] ^ data_in[47] ^ data_in[48] ^ data_in[49] ^ data_in[50] ^ data_in[51] ^ data_in[52] ^ data_in[53] ^ data_in[54] ^ data_in[55] ^ data_in[56] ^ data_in[57] ^ data_in[58] ^ data_in[59] ^ data_in[60] ^ data_in[61] ^ data_in[62] ^ data_in[63] ^ data_in[64] ^ data_in[65] ^ data_in[66] ^ data_in[67] ^ data_in[68] ^ data_in[69] ^ data_in[70] ^ data_in[71] ^ data_in[72] ^ data_in[73] ^ data_in[74] ^ data_in[75] ^ data_in[76] ^ data_in[77] ^ data_in[78] ^ data_in[79] ^ data_in[80] ^ data_in[81] ^ data_in[82] ^ data_in[83] ^ data_in[84] ^ data_in[85] ^ data_in[86] ^ data_in[87] ^ data_in[88] ^ data_in[89] ^ data_in[90] ^ data_in[91] ^ data_in[92] ^ data_in[93] ^ data_in[94] ^ data_in[95] ^ data_in[96] ^ data_in[97] ^ data_in[98] ^ data_in[99] ^ data_in[100] ^ data_in[101] ^ data_in[102] ^ data_in[103] ^ data_in[104] ^ data_in[105] ^ data_in[106] ^ data_in[107] ^ data_in[108] ^ data_in[109] ^ data_in[110] ^ data_in[111] ^ data_in[112] ^ data_in[113] ^ data_in[114] ^ data_in[115] ^ data_in[116] ^ data_in[117] ^ data_in[118] ^ data_in[119] ^ data_in[120] ^ data_in[121] ^ data_in[122] ^ data_in[123] ^ data_in[124] ^ data_in[125] ^ data_in[126] ^ data_in[127] ^ data_in[128] ^ data_in[129] ^ data_in[130] ^ data_in[131] ^ data_in[132] ^ data_in[133] ^ data_in[134] ^ data_in[135] ^ data_in[136] ^ data_in[137] ^ data_in[138] ^ data_in[139] ^ data_in[140] ^ data_in[141] ^ data_in[142] ^ data_in[143] ^ data_in[144] ^ data_in[145] ^ data_in[146] ^ data_in[147] ^ data_in[148] ^ data_in[149] ^ data_in[150] ^ data_in[151] ^ data_in[152] ^ data_in[153] ^ data_in[154] ^ data_in[155] ^ data_in[156] ^ data_in[157] ^ data_in[158] ^ data_in[159] ^ data_in[160] ^ data_in[161] ^ data_in[162] ^ data_in[163] ^ data_in[164] ^ data_in[165] ^ data_in[166] ^ data_in[167] ^ data_in[168] ^ data_in[169] ^ data_in[170] ^ data_in[171] ^ data_in[172] ^ data_in[173] ^ data_in[174] ^ data_in[175] ^ data_in[176] ^ data_in[177] ^ data_in[178] ^ data_in[179] ^ data_in[180] ^ data_in[181] ^ data_in[182] ^ data_in[183] ^ data_in[184] ^ data_in[185] ^ data_in[186] ^ data_in[187] ^ data_in[188] ^ data_in[189] ^ data_in[190] ^ data_in[191] ^ data_in[192] ^ data_in[193] ^ data_in[194] ^ data_in[195] ^ data_in[196] ^ data_in[197] ^ data_in[198] ^ data_in[199] ^ data_in[200] ^ data_in[201] ^ data_in[202] ^ data_in[203] ^ data_in[204] ^ data_in[205] ^ data_in[206] ^ data_in[207] ^ data_in[208] ^ data_in[209] ^ data_in[210] ^ data_in[211] ^ data_in[212] ^ data_in[213] ^ data_in[214] ^ data_in[215] ^ data_in[216] ^ data_in[217] ^ data_in[218] ^ data_in[219] ^ data_in[220] ^ data_in[221] ^ data_in[222] ^ data_in[223] ^ data_in[224] ^ data_in[225] ^ data_in[226] ^ data_in[227] ^ data_in[228] ^ data_in[229] ^ data_in[230] ^ data_in[231] ^ data_in[232] ^ data_in[233] ^ data_in[234] ^ data_in[235] ^ data_in[236] ^ data_in[237] ^ data_in[238] ^ data_in[239] ^ data_in[240] ^ data_in[241] ^ data_in[242] ^ data_in[243] ^ data_in[244] ^ data_in[245] ^ data_in[246] ^ data_in[247] ^ data_in[248] ^ data_in[249] ^ data_in[250] ^ data_in[251] ^ data_in[252] ^ data_in[253] ^ data_in[254] ^ data_in[255] ^ data_in[256] ^ data_in[257] ^ data_in[258] ^ data_in[259] ^ data_in[260] ^ data_in[261] ^ data_in[262] ^ data_in[263] ^ data_in[264] ^ data_in[265] ^ data_in[266] ^ data_in[267] ^ data_in[268] ^ data_in[269] ^ data_in[270] ^ data_in[271] ^ data_in[272] ^ data_in[273] ^ data_in[274] ^ data_in[275] ^ data_in[276] ^ data_in[277] ^ data_in[278] ^ data_in[279] ^ data_in[280] ^ data_in[281] ^ data_in[282] ^ data_in[283] ^ data_in[284] ^ data_in[285] ^ data_in[286] ^ data_in[287] ^ data_in[288] ^ data_in[289] ^ data_in[290] ^ data_in[291] ^ data_in[292] ^ data_in[293] ^ data_in[294] ^ data_in[295] ^ data_in[296] ^ data_in[297] ^ data_in[298] ^ data_in[299] ^ data_in[300] ^ data_in[301] ^ data_in[302] ^ data_in[303] ^ data_in[304] ^ data_in[305] ^ data_in[306] ^ data_in[307] ^ data_in[308] ^ data_in[309] ^ data_in[310] ^ data_in[311] ^ data_in[312] ^ data_in[313] ^ data_in[314] ^ data_in[315] ^ data_in[316] ^ data_in[317] ^ data_in[318] ^ data_in[319] ^ data_in[320] ^ data_in[321] ^ data_in[322] ^ data_in[323] ^ data_in[324] ^ data_in[325] ^ data_in[326] ^ data_in[327] ^ data_in[328] ^ data_in[329] ^ data_in[330] ^ data_in[331] ^ data_in[332] ^ data_in[333] ^ data_in[334] ^ data_in[335] ^ data_in[336] ^ data_in[337] ^ data_in[338] ^ data_in[339] ^ data_in[340] ^ data_in[341] ^ data_in[342] ^ data_in[343] ^ data_in[344] ^ data_in[345] ^ data_in[346] ^ data_in[347] ^ data_in[348] ^ data_in[349] ^ data_in[350] ^ data_in[351] ^ data_in[352] ^ data_in[353] ^ data_in[354] ^ data_in[355] ^ data_in[356] ^ data_in[357] ^ data_in[358] ^ data_in[359] ^ data_in[360] ^ data_in[361] ^ data_in[362] ^ data_in[363] ^ data_in[364] ^ data_in[365] ^ data_in[366] ^ data_in[367] ^ data_in[368] ^ data_in[369] ^ data_in[370] ^ data_in[371] ^ data_in[372] ^ data_in[373] ^ data_in[374] ^ data_in[375] ^ data_in[376] ^ data_in[377] ^ data_in[378] ^ data_in[379] ^ data_in[380] ^ data_in[381] ^ data_in[382] ^ data_in[383] ^ data_in[384] ^ data_in[385] ^ data_in[386] ^ data_in[387] ^ data_in[388] ^ data_in[389] ^ data_in[390] ^ data_in[391] ^ data_in[392] ^ data_in[393] ^ data_in[394] ^ data_in[395] ^ data_in[396] ^ data_in[397] ^ data_in[398] ^ data_in[399] ^ data_in[400] ^ data_in[401] ^ data_in[402] ^ data_in[403] ^ data_in[404] ^ data_in[405] ^ data_in[406] ^ data_in[407] ^ data_in[408] ^ data_in[409] ^ data_in[410] ^ data_in[411] ^ data_in[412] ^ data_in[413] ^ data_in[414] ^ data_in[415] ^ data_in[416] ^ data_in[417] ^ data_in[418] ^ data_in[419] ^ data_in[420] ^ data_in[421] ^ data_in[422] ^ data_in[423] ^ data_in[424] ^ data_in[425] ^ data_in[426] ^ data_in[427] ^ data_in[428] ^ data_in[429] ^ data_in[430] ^ data_in[431] ^ data_in[432] ^ data_in[433] ^ data_in[434] ^ data_in[435] ^ data_in[436] ^ data_in[437] ^ data_in[438] ^ data_in[439] ^ data_in[440] ^ data_in[441] ^ data_in[442] ^ data_in[443] ^ data_in[444] ^ data_in[445] ^ data_in[446] ^ data_in[447] ^ data_in[448] ^ data_in[449] ^ data_in[450] ^ data_in[451] ^ data_in[452] ^ data_in[453] ^ data_in[454] ^ data_in[455] ^ data_in[456] ^ data_in[457] ^ data_in[458] ^ data_in[459] ^ data_in[460] ^ data_in[461] ^ data_in[462] ^ data_in[463] ^ data_in[464] ^ data_in[465] ^ data_in[466] ^ data_in[467] ^ data_in[468] ^ data_in[469] ^ data_in[470] ^ data_in[471] ^ data_in[472] ^ data_in[473] ^ data_in[474] ^ data_in[475] ^ data_in[476] ^ data_in[477] ^ data_in[478] ^ data_in[479] ^ data_in[480] ^ data_in[481] ^ data_in[482] ^ data_in[483] ^ data_in[484] ^ data_in[485] ^ data_in[486] ^ data_in[487] ^ data_in[488] ^ data_in[489] ^ data_in[490] ^ data_in[491] ^ data_in[492] ^ data_in[493] ^ data_in[494] ^ data_in[495] ^ data_in[496] ^ data_in[497] ^ data_in[498] ^ data_in[499] ^ data_in[500] ^ data_in[501] ^ checker_in[0] ^ checker_in[1] ^ checker_in[2] ^ checker_in[3] ^ checker_in[4] ^ checker_in[5] ^ checker_in[6] ^ checker_in[7] ^ checker_in[8] ;

end // always(*)
endmodule


module data_mem_10(clock, reset, we, data_in, data_out);

input              clock;
input              reset;
input              we;
input      [ 501:0] data_in;
output reg [ 501:0] data_out;

always @(posedge clock) begin
    if (reset) begin
        data_out <= 0;
    end
    else if (we) begin
        data_out <= data_in;
    end
end
endmodule


module ecc_mem_10(clock, reset, we, checker_in, parity_in, checker_out, parity_out);

input              clock;
input              reset;
input              we;
input      [  8:0] checker_in;
input              parity_in;
output reg [  8:0] checker_out;
output reg         parity_out;

always @(posedge clock) begin
    if (reset) begin
        checker_out <= 0;
        parity_out <= 0;
    end
    else if (we) begin
        checker_out <= checker_in;
        parity_out <= parity_in;
    end
end
endmodule


module ecc_corrector_10(data_out, checker_out, parity_out, correct_data_out, error);

input      [ 501:0] data_out;
input      [  8:0] checker_out;
input              parity_out;
output reg [ 501:0] correct_data_out;
output reg         error;

reg        [  8:0] syndrome;
reg                parity;

always @(*) begin
    syndrome[0] = data_out[501] ^ data_out[500] ^ data_out[498] ^ data_out[497] ^ data_out[495] ^ data_out[493] ^ data_out[491] ^ data_out[490] ^ data_out[488] ^ data_out[486] ^ data_out[484] ^ data_out[482] ^ data_out[480] ^ data_out[478] ^ data_out[476] ^ data_out[475] ^ data_out[473] ^ data_out[471] ^ data_out[469] ^ data_out[467] ^ data_out[465] ^ data_out[463] ^ data_out[461] ^ data_out[459] ^ data_out[457] ^ data_out[455] ^ data_out[453] ^ data_out[451] ^ data_out[449] ^ data_out[447] ^ data_out[445] ^ data_out[444] ^ data_out[442] ^ data_out[440] ^ data_out[438] ^ data_out[436] ^ data_out[434] ^ data_out[432] ^ data_out[430] ^ data_out[428] ^ data_out[426] ^ data_out[424] ^ data_out[422] ^ data_out[420] ^ data_out[418] ^ data_out[416] ^ data_out[414] ^ data_out[412] ^ data_out[410] ^ data_out[408] ^ data_out[406] ^ data_out[404] ^ data_out[402] ^ data_out[400] ^ data_out[398] ^ data_out[396] ^ data_out[394] ^ data_out[392] ^ data_out[390] ^ data_out[388] ^ data_out[386] ^ data_out[384] ^ data_out[382] ^ data_out[381] ^ data_out[379] ^ data_out[377] ^ data_out[375] ^ data_out[373] ^ data_out[371] ^ data_out[369] ^ data_out[367] ^ data_out[365] ^ data_out[363] ^ data_out[361] ^ data_out[359] ^ data_out[357] ^ data_out[355] ^ data_out[353] ^ data_out[351] ^ data_out[349] ^ data_out[347] ^ data_out[345] ^ data_out[343] ^ data_out[341] ^ data_out[339] ^ data_out[337] ^ data_out[335] ^ data_out[333] ^ data_out[331] ^ data_out[329] ^ data_out[327] ^ data_out[325] ^ data_out[323] ^ data_out[321] ^ data_out[319] ^ data_out[317] ^ data_out[315] ^ data_out[313] ^ data_out[311] ^ data_out[309] ^ data_out[307] ^ data_out[305] ^ data_out[303] ^ data_out[301] ^ data_out[299] ^ data_out[297] ^ data_out[295] ^ data_out[293] ^ data_out[291] ^ data_out[289] ^ data_out[287] ^ data_out[285] ^ data_out[283] ^ data_out[281] ^ data_out[279] ^ data_out[277] ^ data_out[275] ^ data_out[273] ^ data_out[271] ^ data_out[269] ^ data_out[267] ^ data_out[265] ^ data_out[263] ^ data_out[261] ^ data_out[259] ^ data_out[257] ^ data_out[255] ^ data_out[254] ^ data_out[252] ^ data_out[250] ^ data_out[248] ^ data_out[246] ^ data_out[244] ^ data_out[242] ^ data_out[240] ^ data_out[238] ^ data_out[236] ^ data_out[234] ^ data_out[232] ^ data_out[230] ^ data_out[228] ^ data_out[226] ^ data_out[224] ^ data_out[222] ^ data_out[220] ^ data_out[218] ^ data_out[216] ^ data_out[214] ^ data_out[212] ^ data_out[210] ^ data_out[208] ^ data_out[206] ^ data_out[204] ^ data_out[202] ^ data_out[200] ^ data_out[198] ^ data_out[196] ^ data_out[194] ^ data_out[192] ^ data_out[190] ^ data_out[188] ^ data_out[186] ^ data_out[184] ^ data_out[182] ^ data_out[180] ^ data_out[178] ^ data_out[176] ^ data_out[174] ^ data_out[172] ^ data_out[170] ^ data_out[168] ^ data_out[166] ^ data_out[164] ^ data_out[162] ^ data_out[160] ^ data_out[158] ^ data_out[156] ^ data_out[154] ^ data_out[152] ^ data_out[150] ^ data_out[148] ^ data_out[146] ^ data_out[144] ^ data_out[142] ^ data_out[140] ^ data_out[138] ^ data_out[136] ^ data_out[134] ^ data_out[132] ^ data_out[130] ^ data_out[128] ^ data_out[126] ^ data_out[124] ^ data_out[122] ^ data_out[120] ^ data_out[118] ^ data_out[116] ^ data_out[114] ^ data_out[112] ^ data_out[110] ^ data_out[108] ^ data_out[106] ^ data_out[104] ^ data_out[102] ^ data_out[100] ^ data_out[98] ^ data_out[96] ^ data_out[94] ^ data_out[92] ^ data_out[90] ^ data_out[88] ^ data_out[86] ^ data_out[84] ^ data_out[82] ^ data_out[80] ^ data_out[78] ^ data_out[76] ^ data_out[74] ^ data_out[72] ^ data_out[70] ^ data_out[68] ^ data_out[66] ^ data_out[64] ^ data_out[62] ^ data_out[60] ^ data_out[58] ^ data_out[56] ^ data_out[54] ^ data_out[52] ^ data_out[50] ^ data_out[48] ^ data_out[46] ^ data_out[44] ^ data_out[42] ^ data_out[40] ^ data_out[38] ^ data_out[36] ^ data_out[34] ^ data_out[32] ^ data_out[30] ^ data_out[28] ^ data_out[26] ^ data_out[24] ^ data_out[22] ^ data_out[20] ^ data_out[18] ^ data_out[16] ^ data_out[14] ^ data_out[12] ^ data_out[10] ^ data_out[8] ^ data_out[6] ^ data_out[4] ^ data_out[2] ^ data_out[0] ^ checker_out[0] ;
    syndrome[1] = data_out[501] ^ data_out[499] ^ data_out[498] ^ data_out[496] ^ data_out[495] ^ data_out[492] ^ data_out[491] ^ data_out[489] ^ data_out[488] ^ data_out[485] ^ data_out[484] ^ data_out[481] ^ data_out[480] ^ data_out[477] ^ data_out[476] ^ data_out[474] ^ data_out[473] ^ data_out[470] ^ data_out[469] ^ data_out[466] ^ data_out[465] ^ data_out[462] ^ data_out[461] ^ data_out[458] ^ data_out[457] ^ data_out[454] ^ data_out[453] ^ data_out[450] ^ data_out[449] ^ data_out[446] ^ data_out[445] ^ data_out[443] ^ data_out[442] ^ data_out[439] ^ data_out[438] ^ data_out[435] ^ data_out[434] ^ data_out[431] ^ data_out[430] ^ data_out[427] ^ data_out[426] ^ data_out[423] ^ data_out[422] ^ data_out[419] ^ data_out[418] ^ data_out[415] ^ data_out[414] ^ data_out[411] ^ data_out[410] ^ data_out[407] ^ data_out[406] ^ data_out[403] ^ data_out[402] ^ data_out[399] ^ data_out[398] ^ data_out[395] ^ data_out[394] ^ data_out[391] ^ data_out[390] ^ data_out[387] ^ data_out[386] ^ data_out[383] ^ data_out[382] ^ data_out[380] ^ data_out[379] ^ data_out[376] ^ data_out[375] ^ data_out[372] ^ data_out[371] ^ data_out[368] ^ data_out[367] ^ data_out[364] ^ data_out[363] ^ data_out[360] ^ data_out[359] ^ data_out[356] ^ data_out[355] ^ data_out[352] ^ data_out[351] ^ data_out[348] ^ data_out[347] ^ data_out[344] ^ data_out[343] ^ data_out[340] ^ data_out[339] ^ data_out[336] ^ data_out[335] ^ data_out[332] ^ data_out[331] ^ data_out[328] ^ data_out[327] ^ data_out[324] ^ data_out[323] ^ data_out[320] ^ data_out[319] ^ data_out[316] ^ data_out[315] ^ data_out[312] ^ data_out[311] ^ data_out[308] ^ data_out[307] ^ data_out[304] ^ data_out[303] ^ data_out[300] ^ data_out[299] ^ data_out[296] ^ data_out[295] ^ data_out[292] ^ data_out[291] ^ data_out[288] ^ data_out[287] ^ data_out[284] ^ data_out[283] ^ data_out[280] ^ data_out[279] ^ data_out[276] ^ data_out[275] ^ data_out[272] ^ data_out[271] ^ data_out[268] ^ data_out[267] ^ data_out[264] ^ data_out[263] ^ data_out[260] ^ data_out[259] ^ data_out[256] ^ data_out[255] ^ data_out[253] ^ data_out[252] ^ data_out[249] ^ data_out[248] ^ data_out[245] ^ data_out[244] ^ data_out[241] ^ data_out[240] ^ data_out[237] ^ data_out[236] ^ data_out[233] ^ data_out[232] ^ data_out[229] ^ data_out[228] ^ data_out[225] ^ data_out[224] ^ data_out[221] ^ data_out[220] ^ data_out[217] ^ data_out[216] ^ data_out[213] ^ data_out[212] ^ data_out[209] ^ data_out[208] ^ data_out[205] ^ data_out[204] ^ data_out[201] ^ data_out[200] ^ data_out[197] ^ data_out[196] ^ data_out[193] ^ data_out[192] ^ data_out[189] ^ data_out[188] ^ data_out[185] ^ data_out[184] ^ data_out[181] ^ data_out[180] ^ data_out[177] ^ data_out[176] ^ data_out[173] ^ data_out[172] ^ data_out[169] ^ data_out[168] ^ data_out[165] ^ data_out[164] ^ data_out[161] ^ data_out[160] ^ data_out[157] ^ data_out[156] ^ data_out[153] ^ data_out[152] ^ data_out[149] ^ data_out[148] ^ data_out[145] ^ data_out[144] ^ data_out[141] ^ data_out[140] ^ data_out[137] ^ data_out[136] ^ data_out[133] ^ data_out[132] ^ data_out[129] ^ data_out[128] ^ data_out[125] ^ data_out[124] ^ data_out[121] ^ data_out[120] ^ data_out[117] ^ data_out[116] ^ data_out[113] ^ data_out[112] ^ data_out[109] ^ data_out[108] ^ data_out[105] ^ data_out[104] ^ data_out[101] ^ data_out[100] ^ data_out[97] ^ data_out[96] ^ data_out[93] ^ data_out[92] ^ data_out[89] ^ data_out[88] ^ data_out[85] ^ data_out[84] ^ data_out[81] ^ data_out[80] ^ data_out[77] ^ data_out[76] ^ data_out[73] ^ data_out[72] ^ data_out[69] ^ data_out[68] ^ data_out[65] ^ data_out[64] ^ data_out[61] ^ data_out[60] ^ data_out[57] ^ data_out[56] ^ data_out[53] ^ data_out[52] ^ data_out[49] ^ data_out[48] ^ data_out[45] ^ data_out[44] ^ data_out[41] ^ data_out[40] ^ data_out[37] ^ data_out[36] ^ data_out[33] ^ data_out[32] ^ data_out[29] ^ data_out[28] ^ data_out[25] ^ data_out[24] ^ data_out[21] ^ data_out[20] ^ data_out[17] ^ data_out[16] ^ data_out[13] ^ data_out[12] ^ data_out[9] ^ data_out[8] ^ data_out[5] ^ data_out[4] ^ data_out[1] ^ data_out[0] ^ checker_out[1] ;
    syndrome[2] = data_out[500] ^ data_out[499] ^ data_out[498] ^ data_out[494] ^ data_out[493] ^ data_out[492] ^ data_out[491] ^ data_out[487] ^ data_out[486] ^ data_out[485] ^ data_out[484] ^ data_out[479] ^ data_out[478] ^ data_out[477] ^ data_out[476] ^ data_out[472] ^ data_out[471] ^ data_out[470] ^ data_out[469] ^ data_out[464] ^ data_out[463] ^ data_out[462] ^ data_out[461] ^ data_out[456] ^ data_out[455] ^ data_out[454] ^ data_out[453] ^ data_out[448] ^ data_out[447] ^ data_out[446] ^ data_out[445] ^ data_out[441] ^ data_out[440] ^ data_out[439] ^ data_out[438] ^ data_out[433] ^ data_out[432] ^ data_out[431] ^ data_out[430] ^ data_out[425] ^ data_out[424] ^ data_out[423] ^ data_out[422] ^ data_out[417] ^ data_out[416] ^ data_out[415] ^ data_out[414] ^ data_out[409] ^ data_out[408] ^ data_out[407] ^ data_out[406] ^ data_out[401] ^ data_out[400] ^ data_out[399] ^ data_out[398] ^ data_out[393] ^ data_out[392] ^ data_out[391] ^ data_out[390] ^ data_out[385] ^ data_out[384] ^ data_out[383] ^ data_out[382] ^ data_out[378] ^ data_out[377] ^ data_out[376] ^ data_out[375] ^ data_out[370] ^ data_out[369] ^ data_out[368] ^ data_out[367] ^ data_out[362] ^ data_out[361] ^ data_out[360] ^ data_out[359] ^ data_out[354] ^ data_out[353] ^ data_out[352] ^ data_out[351] ^ data_out[346] ^ data_out[345] ^ data_out[344] ^ data_out[343] ^ data_out[338] ^ data_out[337] ^ data_out[336] ^ data_out[335] ^ data_out[330] ^ data_out[329] ^ data_out[328] ^ data_out[327] ^ data_out[322] ^ data_out[321] ^ data_out[320] ^ data_out[319] ^ data_out[314] ^ data_out[313] ^ data_out[312] ^ data_out[311] ^ data_out[306] ^ data_out[305] ^ data_out[304] ^ data_out[303] ^ data_out[298] ^ data_out[297] ^ data_out[296] ^ data_out[295] ^ data_out[290] ^ data_out[289] ^ data_out[288] ^ data_out[287] ^ data_out[282] ^ data_out[281] ^ data_out[280] ^ data_out[279] ^ data_out[274] ^ data_out[273] ^ data_out[272] ^ data_out[271] ^ data_out[266] ^ data_out[265] ^ data_out[264] ^ data_out[263] ^ data_out[258] ^ data_out[257] ^ data_out[256] ^ data_out[255] ^ data_out[251] ^ data_out[250] ^ data_out[249] ^ data_out[248] ^ data_out[243] ^ data_out[242] ^ data_out[241] ^ data_out[240] ^ data_out[235] ^ data_out[234] ^ data_out[233] ^ data_out[232] ^ data_out[227] ^ data_out[226] ^ data_out[225] ^ data_out[224] ^ data_out[219] ^ data_out[218] ^ data_out[217] ^ data_out[216] ^ data_out[211] ^ data_out[210] ^ data_out[209] ^ data_out[208] ^ data_out[203] ^ data_out[202] ^ data_out[201] ^ data_out[200] ^ data_out[195] ^ data_out[194] ^ data_out[193] ^ data_out[192] ^ data_out[187] ^ data_out[186] ^ data_out[185] ^ data_out[184] ^ data_out[179] ^ data_out[178] ^ data_out[177] ^ data_out[176] ^ data_out[171] ^ data_out[170] ^ data_out[169] ^ data_out[168] ^ data_out[163] ^ data_out[162] ^ data_out[161] ^ data_out[160] ^ data_out[155] ^ data_out[154] ^ data_out[153] ^ data_out[152] ^ data_out[147] ^ data_out[146] ^ data_out[145] ^ data_out[144] ^ data_out[139] ^ data_out[138] ^ data_out[137] ^ data_out[136] ^ data_out[131] ^ data_out[130] ^ data_out[129] ^ data_out[128] ^ data_out[123] ^ data_out[122] ^ data_out[121] ^ data_out[120] ^ data_out[115] ^ data_out[114] ^ data_out[113] ^ data_out[112] ^ data_out[107] ^ data_out[106] ^ data_out[105] ^ data_out[104] ^ data_out[99] ^ data_out[98] ^ data_out[97] ^ data_out[96] ^ data_out[91] ^ data_out[90] ^ data_out[89] ^ data_out[88] ^ data_out[83] ^ data_out[82] ^ data_out[81] ^ data_out[80] ^ data_out[75] ^ data_out[74] ^ data_out[73] ^ data_out[72] ^ data_out[67] ^ data_out[66] ^ data_out[65] ^ data_out[64] ^ data_out[59] ^ data_out[58] ^ data_out[57] ^ data_out[56] ^ data_out[51] ^ data_out[50] ^ data_out[49] ^ data_out[48] ^ data_out[43] ^ data_out[42] ^ data_out[41] ^ data_out[40] ^ data_out[35] ^ data_out[34] ^ data_out[33] ^ data_out[32] ^ data_out[27] ^ data_out[26] ^ data_out[25] ^ data_out[24] ^ data_out[19] ^ data_out[18] ^ data_out[17] ^ data_out[16] ^ data_out[11] ^ data_out[10] ^ data_out[9] ^ data_out[8] ^ data_out[3] ^ data_out[2] ^ data_out[1] ^ data_out[0] ^ checker_out[2] ;
    syndrome[3] = data_out[497] ^ data_out[496] ^ data_out[495] ^ data_out[494] ^ data_out[493] ^ data_out[492] ^ data_out[491] ^ data_out[483] ^ data_out[482] ^ data_out[481] ^ data_out[480] ^ data_out[479] ^ data_out[478] ^ data_out[477] ^ data_out[476] ^ data_out[468] ^ data_out[467] ^ data_out[466] ^ data_out[465] ^ data_out[464] ^ data_out[463] ^ data_out[462] ^ data_out[461] ^ data_out[452] ^ data_out[451] ^ data_out[450] ^ data_out[449] ^ data_out[448] ^ data_out[447] ^ data_out[446] ^ data_out[445] ^ data_out[437] ^ data_out[436] ^ data_out[435] ^ data_out[434] ^ data_out[433] ^ data_out[432] ^ data_out[431] ^ data_out[430] ^ data_out[421] ^ data_out[420] ^ data_out[419] ^ data_out[418] ^ data_out[417] ^ data_out[416] ^ data_out[415] ^ data_out[414] ^ data_out[405] ^ data_out[404] ^ data_out[403] ^ data_out[402] ^ data_out[401] ^ data_out[400] ^ data_out[399] ^ data_out[398] ^ data_out[389] ^ data_out[388] ^ data_out[387] ^ data_out[386] ^ data_out[385] ^ data_out[384] ^ data_out[383] ^ data_out[382] ^ data_out[374] ^ data_out[373] ^ data_out[372] ^ data_out[371] ^ data_out[370] ^ data_out[369] ^ data_out[368] ^ data_out[367] ^ data_out[358] ^ data_out[357] ^ data_out[356] ^ data_out[355] ^ data_out[354] ^ data_out[353] ^ data_out[352] ^ data_out[351] ^ data_out[342] ^ data_out[341] ^ data_out[340] ^ data_out[339] ^ data_out[338] ^ data_out[337] ^ data_out[336] ^ data_out[335] ^ data_out[326] ^ data_out[325] ^ data_out[324] ^ data_out[323] ^ data_out[322] ^ data_out[321] ^ data_out[320] ^ data_out[319] ^ data_out[310] ^ data_out[309] ^ data_out[308] ^ data_out[307] ^ data_out[306] ^ data_out[305] ^ data_out[304] ^ data_out[303] ^ data_out[294] ^ data_out[293] ^ data_out[292] ^ data_out[291] ^ data_out[290] ^ data_out[289] ^ data_out[288] ^ data_out[287] ^ data_out[278] ^ data_out[277] ^ data_out[276] ^ data_out[275] ^ data_out[274] ^ data_out[273] ^ data_out[272] ^ data_out[271] ^ data_out[262] ^ data_out[261] ^ data_out[260] ^ data_out[259] ^ data_out[258] ^ data_out[257] ^ data_out[256] ^ data_out[255] ^ data_out[247] ^ data_out[246] ^ data_out[245] ^ data_out[244] ^ data_out[243] ^ data_out[242] ^ data_out[241] ^ data_out[240] ^ data_out[231] ^ data_out[230] ^ data_out[229] ^ data_out[228] ^ data_out[227] ^ data_out[226] ^ data_out[225] ^ data_out[224] ^ data_out[215] ^ data_out[214] ^ data_out[213] ^ data_out[212] ^ data_out[211] ^ data_out[210] ^ data_out[209] ^ data_out[208] ^ data_out[199] ^ data_out[198] ^ data_out[197] ^ data_out[196] ^ data_out[195] ^ data_out[194] ^ data_out[193] ^ data_out[192] ^ data_out[183] ^ data_out[182] ^ data_out[181] ^ data_out[180] ^ data_out[179] ^ data_out[178] ^ data_out[177] ^ data_out[176] ^ data_out[167] ^ data_out[166] ^ data_out[165] ^ data_out[164] ^ data_out[163] ^ data_out[162] ^ data_out[161] ^ data_out[160] ^ data_out[151] ^ data_out[150] ^ data_out[149] ^ data_out[148] ^ data_out[147] ^ data_out[146] ^ data_out[145] ^ data_out[144] ^ data_out[135] ^ data_out[134] ^ data_out[133] ^ data_out[132] ^ data_out[131] ^ data_out[130] ^ data_out[129] ^ data_out[128] ^ data_out[119] ^ data_out[118] ^ data_out[117] ^ data_out[116] ^ data_out[115] ^ data_out[114] ^ data_out[113] ^ data_out[112] ^ data_out[103] ^ data_out[102] ^ data_out[101] ^ data_out[100] ^ data_out[99] ^ data_out[98] ^ data_out[97] ^ data_out[96] ^ data_out[87] ^ data_out[86] ^ data_out[85] ^ data_out[84] ^ data_out[83] ^ data_out[82] ^ data_out[81] ^ data_out[80] ^ data_out[71] ^ data_out[70] ^ data_out[69] ^ data_out[68] ^ data_out[67] ^ data_out[66] ^ data_out[65] ^ data_out[64] ^ data_out[55] ^ data_out[54] ^ data_out[53] ^ data_out[52] ^ data_out[51] ^ data_out[50] ^ data_out[49] ^ data_out[48] ^ data_out[39] ^ data_out[38] ^ data_out[37] ^ data_out[36] ^ data_out[35] ^ data_out[34] ^ data_out[33] ^ data_out[32] ^ data_out[23] ^ data_out[22] ^ data_out[21] ^ data_out[20] ^ data_out[19] ^ data_out[18] ^ data_out[17] ^ data_out[16] ^ data_out[7] ^ data_out[6] ^ data_out[5] ^ data_out[4] ^ data_out[3] ^ data_out[2] ^ data_out[1] ^ data_out[0] ^ checker_out[3] ;
    syndrome[4] = data_out[490] ^ data_out[489] ^ data_out[488] ^ data_out[487] ^ data_out[486] ^ data_out[485] ^ data_out[484] ^ data_out[483] ^ data_out[482] ^ data_out[481] ^ data_out[480] ^ data_out[479] ^ data_out[478] ^ data_out[477] ^ data_out[476] ^ data_out[460] ^ data_out[459] ^ data_out[458] ^ data_out[457] ^ data_out[456] ^ data_out[455] ^ data_out[454] ^ data_out[453] ^ data_out[452] ^ data_out[451] ^ data_out[450] ^ data_out[449] ^ data_out[448] ^ data_out[447] ^ data_out[446] ^ data_out[445] ^ data_out[429] ^ data_out[428] ^ data_out[427] ^ data_out[426] ^ data_out[425] ^ data_out[424] ^ data_out[423] ^ data_out[422] ^ data_out[421] ^ data_out[420] ^ data_out[419] ^ data_out[418] ^ data_out[417] ^ data_out[416] ^ data_out[415] ^ data_out[414] ^ data_out[397] ^ data_out[396] ^ data_out[395] ^ data_out[394] ^ data_out[393] ^ data_out[392] ^ data_out[391] ^ data_out[390] ^ data_out[389] ^ data_out[388] ^ data_out[387] ^ data_out[386] ^ data_out[385] ^ data_out[384] ^ data_out[383] ^ data_out[382] ^ data_out[366] ^ data_out[365] ^ data_out[364] ^ data_out[363] ^ data_out[362] ^ data_out[361] ^ data_out[360] ^ data_out[359] ^ data_out[358] ^ data_out[357] ^ data_out[356] ^ data_out[355] ^ data_out[354] ^ data_out[353] ^ data_out[352] ^ data_out[351] ^ data_out[334] ^ data_out[333] ^ data_out[332] ^ data_out[331] ^ data_out[330] ^ data_out[329] ^ data_out[328] ^ data_out[327] ^ data_out[326] ^ data_out[325] ^ data_out[324] ^ data_out[323] ^ data_out[322] ^ data_out[321] ^ data_out[320] ^ data_out[319] ^ data_out[302] ^ data_out[301] ^ data_out[300] ^ data_out[299] ^ data_out[298] ^ data_out[297] ^ data_out[296] ^ data_out[295] ^ data_out[294] ^ data_out[293] ^ data_out[292] ^ data_out[291] ^ data_out[290] ^ data_out[289] ^ data_out[288] ^ data_out[287] ^ data_out[270] ^ data_out[269] ^ data_out[268] ^ data_out[267] ^ data_out[266] ^ data_out[265] ^ data_out[264] ^ data_out[263] ^ data_out[262] ^ data_out[261] ^ data_out[260] ^ data_out[259] ^ data_out[258] ^ data_out[257] ^ data_out[256] ^ data_out[255] ^ data_out[239] ^ data_out[238] ^ data_out[237] ^ data_out[236] ^ data_out[235] ^ data_out[234] ^ data_out[233] ^ data_out[232] ^ data_out[231] ^ data_out[230] ^ data_out[229] ^ data_out[228] ^ data_out[227] ^ data_out[226] ^ data_out[225] ^ data_out[224] ^ data_out[207] ^ data_out[206] ^ data_out[205] ^ data_out[204] ^ data_out[203] ^ data_out[202] ^ data_out[201] ^ data_out[200] ^ data_out[199] ^ data_out[198] ^ data_out[197] ^ data_out[196] ^ data_out[195] ^ data_out[194] ^ data_out[193] ^ data_out[192] ^ data_out[175] ^ data_out[174] ^ data_out[173] ^ data_out[172] ^ data_out[171] ^ data_out[170] ^ data_out[169] ^ data_out[168] ^ data_out[167] ^ data_out[166] ^ data_out[165] ^ data_out[164] ^ data_out[163] ^ data_out[162] ^ data_out[161] ^ data_out[160] ^ data_out[143] ^ data_out[142] ^ data_out[141] ^ data_out[140] ^ data_out[139] ^ data_out[138] ^ data_out[137] ^ data_out[136] ^ data_out[135] ^ data_out[134] ^ data_out[133] ^ data_out[132] ^ data_out[131] ^ data_out[130] ^ data_out[129] ^ data_out[128] ^ data_out[111] ^ data_out[110] ^ data_out[109] ^ data_out[108] ^ data_out[107] ^ data_out[106] ^ data_out[105] ^ data_out[104] ^ data_out[103] ^ data_out[102] ^ data_out[101] ^ data_out[100] ^ data_out[99] ^ data_out[98] ^ data_out[97] ^ data_out[96] ^ data_out[79] ^ data_out[78] ^ data_out[77] ^ data_out[76] ^ data_out[75] ^ data_out[74] ^ data_out[73] ^ data_out[72] ^ data_out[71] ^ data_out[70] ^ data_out[69] ^ data_out[68] ^ data_out[67] ^ data_out[66] ^ data_out[65] ^ data_out[64] ^ data_out[47] ^ data_out[46] ^ data_out[45] ^ data_out[44] ^ data_out[43] ^ data_out[42] ^ data_out[41] ^ data_out[40] ^ data_out[39] ^ data_out[38] ^ data_out[37] ^ data_out[36] ^ data_out[35] ^ data_out[34] ^ data_out[33] ^ data_out[32] ^ data_out[15] ^ data_out[14] ^ data_out[13] ^ data_out[12] ^ data_out[11] ^ data_out[10] ^ data_out[9] ^ data_out[8] ^ data_out[7] ^ data_out[6] ^ data_out[5] ^ data_out[4] ^ data_out[3] ^ data_out[2] ^ data_out[1] ^ data_out[0] ^ checker_out[4] ;
    syndrome[5] = data_out[475] ^ data_out[474] ^ data_out[473] ^ data_out[472] ^ data_out[471] ^ data_out[470] ^ data_out[469] ^ data_out[468] ^ data_out[467] ^ data_out[466] ^ data_out[465] ^ data_out[464] ^ data_out[463] ^ data_out[462] ^ data_out[461] ^ data_out[460] ^ data_out[459] ^ data_out[458] ^ data_out[457] ^ data_out[456] ^ data_out[455] ^ data_out[454] ^ data_out[453] ^ data_out[452] ^ data_out[451] ^ data_out[450] ^ data_out[449] ^ data_out[448] ^ data_out[447] ^ data_out[446] ^ data_out[445] ^ data_out[413] ^ data_out[412] ^ data_out[411] ^ data_out[410] ^ data_out[409] ^ data_out[408] ^ data_out[407] ^ data_out[406] ^ data_out[405] ^ data_out[404] ^ data_out[403] ^ data_out[402] ^ data_out[401] ^ data_out[400] ^ data_out[399] ^ data_out[398] ^ data_out[397] ^ data_out[396] ^ data_out[395] ^ data_out[394] ^ data_out[393] ^ data_out[392] ^ data_out[391] ^ data_out[390] ^ data_out[389] ^ data_out[388] ^ data_out[387] ^ data_out[386] ^ data_out[385] ^ data_out[384] ^ data_out[383] ^ data_out[382] ^ data_out[350] ^ data_out[349] ^ data_out[348] ^ data_out[347] ^ data_out[346] ^ data_out[345] ^ data_out[344] ^ data_out[343] ^ data_out[342] ^ data_out[341] ^ data_out[340] ^ data_out[339] ^ data_out[338] ^ data_out[337] ^ data_out[336] ^ data_out[335] ^ data_out[334] ^ data_out[333] ^ data_out[332] ^ data_out[331] ^ data_out[330] ^ data_out[329] ^ data_out[328] ^ data_out[327] ^ data_out[326] ^ data_out[325] ^ data_out[324] ^ data_out[323] ^ data_out[322] ^ data_out[321] ^ data_out[320] ^ data_out[319] ^ data_out[286] ^ data_out[285] ^ data_out[284] ^ data_out[283] ^ data_out[282] ^ data_out[281] ^ data_out[280] ^ data_out[279] ^ data_out[278] ^ data_out[277] ^ data_out[276] ^ data_out[275] ^ data_out[274] ^ data_out[273] ^ data_out[272] ^ data_out[271] ^ data_out[270] ^ data_out[269] ^ data_out[268] ^ data_out[267] ^ data_out[266] ^ data_out[265] ^ data_out[264] ^ data_out[263] ^ data_out[262] ^ data_out[261] ^ data_out[260] ^ data_out[259] ^ data_out[258] ^ data_out[257] ^ data_out[256] ^ data_out[255] ^ data_out[223] ^ data_out[222] ^ data_out[221] ^ data_out[220] ^ data_out[219] ^ data_out[218] ^ data_out[217] ^ data_out[216] ^ data_out[215] ^ data_out[214] ^ data_out[213] ^ data_out[212] ^ data_out[211] ^ data_out[210] ^ data_out[209] ^ data_out[208] ^ data_out[207] ^ data_out[206] ^ data_out[205] ^ data_out[204] ^ data_out[203] ^ data_out[202] ^ data_out[201] ^ data_out[200] ^ data_out[199] ^ data_out[198] ^ data_out[197] ^ data_out[196] ^ data_out[195] ^ data_out[194] ^ data_out[193] ^ data_out[192] ^ data_out[159] ^ data_out[158] ^ data_out[157] ^ data_out[156] ^ data_out[155] ^ data_out[154] ^ data_out[153] ^ data_out[152] ^ data_out[151] ^ data_out[150] ^ data_out[149] ^ data_out[148] ^ data_out[147] ^ data_out[146] ^ data_out[145] ^ data_out[144] ^ data_out[143] ^ data_out[142] ^ data_out[141] ^ data_out[140] ^ data_out[139] ^ data_out[138] ^ data_out[137] ^ data_out[136] ^ data_out[135] ^ data_out[134] ^ data_out[133] ^ data_out[132] ^ data_out[131] ^ data_out[130] ^ data_out[129] ^ data_out[128] ^ data_out[95] ^ data_out[94] ^ data_out[93] ^ data_out[92] ^ data_out[91] ^ data_out[90] ^ data_out[89] ^ data_out[88] ^ data_out[87] ^ data_out[86] ^ data_out[85] ^ data_out[84] ^ data_out[83] ^ data_out[82] ^ data_out[81] ^ data_out[80] ^ data_out[79] ^ data_out[78] ^ data_out[77] ^ data_out[76] ^ data_out[75] ^ data_out[74] ^ data_out[73] ^ data_out[72] ^ data_out[71] ^ data_out[70] ^ data_out[69] ^ data_out[68] ^ data_out[67] ^ data_out[66] ^ data_out[65] ^ data_out[64] ^ data_out[31] ^ data_out[30] ^ data_out[29] ^ data_out[28] ^ data_out[27] ^ data_out[26] ^ data_out[25] ^ data_out[24] ^ data_out[23] ^ data_out[22] ^ data_out[21] ^ data_out[20] ^ data_out[19] ^ data_out[18] ^ data_out[17] ^ data_out[16] ^ data_out[15] ^ data_out[14] ^ data_out[13] ^ data_out[12] ^ data_out[11] ^ data_out[10] ^ data_out[9] ^ data_out[8] ^ data_out[7] ^ data_out[6] ^ data_out[5] ^ data_out[4] ^ data_out[3] ^ data_out[2] ^ data_out[1] ^ data_out[0] ^ checker_out[5] ;
    syndrome[6] = data_out[444] ^ data_out[443] ^ data_out[442] ^ data_out[441] ^ data_out[440] ^ data_out[439] ^ data_out[438] ^ data_out[437] ^ data_out[436] ^ data_out[435] ^ data_out[434] ^ data_out[433] ^ data_out[432] ^ data_out[431] ^ data_out[430] ^ data_out[429] ^ data_out[428] ^ data_out[427] ^ data_out[426] ^ data_out[425] ^ data_out[424] ^ data_out[423] ^ data_out[422] ^ data_out[421] ^ data_out[420] ^ data_out[419] ^ data_out[418] ^ data_out[417] ^ data_out[416] ^ data_out[415] ^ data_out[414] ^ data_out[413] ^ data_out[412] ^ data_out[411] ^ data_out[410] ^ data_out[409] ^ data_out[408] ^ data_out[407] ^ data_out[406] ^ data_out[405] ^ data_out[404] ^ data_out[403] ^ data_out[402] ^ data_out[401] ^ data_out[400] ^ data_out[399] ^ data_out[398] ^ data_out[397] ^ data_out[396] ^ data_out[395] ^ data_out[394] ^ data_out[393] ^ data_out[392] ^ data_out[391] ^ data_out[390] ^ data_out[389] ^ data_out[388] ^ data_out[387] ^ data_out[386] ^ data_out[385] ^ data_out[384] ^ data_out[383] ^ data_out[382] ^ data_out[318] ^ data_out[317] ^ data_out[316] ^ data_out[315] ^ data_out[314] ^ data_out[313] ^ data_out[312] ^ data_out[311] ^ data_out[310] ^ data_out[309] ^ data_out[308] ^ data_out[307] ^ data_out[306] ^ data_out[305] ^ data_out[304] ^ data_out[303] ^ data_out[302] ^ data_out[301] ^ data_out[300] ^ data_out[299] ^ data_out[298] ^ data_out[297] ^ data_out[296] ^ data_out[295] ^ data_out[294] ^ data_out[293] ^ data_out[292] ^ data_out[291] ^ data_out[290] ^ data_out[289] ^ data_out[288] ^ data_out[287] ^ data_out[286] ^ data_out[285] ^ data_out[284] ^ data_out[283] ^ data_out[282] ^ data_out[281] ^ data_out[280] ^ data_out[279] ^ data_out[278] ^ data_out[277] ^ data_out[276] ^ data_out[275] ^ data_out[274] ^ data_out[273] ^ data_out[272] ^ data_out[271] ^ data_out[270] ^ data_out[269] ^ data_out[268] ^ data_out[267] ^ data_out[266] ^ data_out[265] ^ data_out[264] ^ data_out[263] ^ data_out[262] ^ data_out[261] ^ data_out[260] ^ data_out[259] ^ data_out[258] ^ data_out[257] ^ data_out[256] ^ data_out[255] ^ data_out[191] ^ data_out[190] ^ data_out[189] ^ data_out[188] ^ data_out[187] ^ data_out[186] ^ data_out[185] ^ data_out[184] ^ data_out[183] ^ data_out[182] ^ data_out[181] ^ data_out[180] ^ data_out[179] ^ data_out[178] ^ data_out[177] ^ data_out[176] ^ data_out[175] ^ data_out[174] ^ data_out[173] ^ data_out[172] ^ data_out[171] ^ data_out[170] ^ data_out[169] ^ data_out[168] ^ data_out[167] ^ data_out[166] ^ data_out[165] ^ data_out[164] ^ data_out[163] ^ data_out[162] ^ data_out[161] ^ data_out[160] ^ data_out[159] ^ data_out[158] ^ data_out[157] ^ data_out[156] ^ data_out[155] ^ data_out[154] ^ data_out[153] ^ data_out[152] ^ data_out[151] ^ data_out[150] ^ data_out[149] ^ data_out[148] ^ data_out[147] ^ data_out[146] ^ data_out[145] ^ data_out[144] ^ data_out[143] ^ data_out[142] ^ data_out[141] ^ data_out[140] ^ data_out[139] ^ data_out[138] ^ data_out[137] ^ data_out[136] ^ data_out[135] ^ data_out[134] ^ data_out[133] ^ data_out[132] ^ data_out[131] ^ data_out[130] ^ data_out[129] ^ data_out[128] ^ data_out[63] ^ data_out[62] ^ data_out[61] ^ data_out[60] ^ data_out[59] ^ data_out[58] ^ data_out[57] ^ data_out[56] ^ data_out[55] ^ data_out[54] ^ data_out[53] ^ data_out[52] ^ data_out[51] ^ data_out[50] ^ data_out[49] ^ data_out[48] ^ data_out[47] ^ data_out[46] ^ data_out[45] ^ data_out[44] ^ data_out[43] ^ data_out[42] ^ data_out[41] ^ data_out[40] ^ data_out[39] ^ data_out[38] ^ data_out[37] ^ data_out[36] ^ data_out[35] ^ data_out[34] ^ data_out[33] ^ data_out[32] ^ data_out[31] ^ data_out[30] ^ data_out[29] ^ data_out[28] ^ data_out[27] ^ data_out[26] ^ data_out[25] ^ data_out[24] ^ data_out[23] ^ data_out[22] ^ data_out[21] ^ data_out[20] ^ data_out[19] ^ data_out[18] ^ data_out[17] ^ data_out[16] ^ data_out[15] ^ data_out[14] ^ data_out[13] ^ data_out[12] ^ data_out[11] ^ data_out[10] ^ data_out[9] ^ data_out[8] ^ data_out[7] ^ data_out[6] ^ data_out[5] ^ data_out[4] ^ data_out[3] ^ data_out[2] ^ data_out[1] ^ data_out[0] ^ checker_out[6] ;
    syndrome[7] = data_out[381] ^ data_out[380] ^ data_out[379] ^ data_out[378] ^ data_out[377] ^ data_out[376] ^ data_out[375] ^ data_out[374] ^ data_out[373] ^ data_out[372] ^ data_out[371] ^ data_out[370] ^ data_out[369] ^ data_out[368] ^ data_out[367] ^ data_out[366] ^ data_out[365] ^ data_out[364] ^ data_out[363] ^ data_out[362] ^ data_out[361] ^ data_out[360] ^ data_out[359] ^ data_out[358] ^ data_out[357] ^ data_out[356] ^ data_out[355] ^ data_out[354] ^ data_out[353] ^ data_out[352] ^ data_out[351] ^ data_out[350] ^ data_out[349] ^ data_out[348] ^ data_out[347] ^ data_out[346] ^ data_out[345] ^ data_out[344] ^ data_out[343] ^ data_out[342] ^ data_out[341] ^ data_out[340] ^ data_out[339] ^ data_out[338] ^ data_out[337] ^ data_out[336] ^ data_out[335] ^ data_out[334] ^ data_out[333] ^ data_out[332] ^ data_out[331] ^ data_out[330] ^ data_out[329] ^ data_out[328] ^ data_out[327] ^ data_out[326] ^ data_out[325] ^ data_out[324] ^ data_out[323] ^ data_out[322] ^ data_out[321] ^ data_out[320] ^ data_out[319] ^ data_out[318] ^ data_out[317] ^ data_out[316] ^ data_out[315] ^ data_out[314] ^ data_out[313] ^ data_out[312] ^ data_out[311] ^ data_out[310] ^ data_out[309] ^ data_out[308] ^ data_out[307] ^ data_out[306] ^ data_out[305] ^ data_out[304] ^ data_out[303] ^ data_out[302] ^ data_out[301] ^ data_out[300] ^ data_out[299] ^ data_out[298] ^ data_out[297] ^ data_out[296] ^ data_out[295] ^ data_out[294] ^ data_out[293] ^ data_out[292] ^ data_out[291] ^ data_out[290] ^ data_out[289] ^ data_out[288] ^ data_out[287] ^ data_out[286] ^ data_out[285] ^ data_out[284] ^ data_out[283] ^ data_out[282] ^ data_out[281] ^ data_out[280] ^ data_out[279] ^ data_out[278] ^ data_out[277] ^ data_out[276] ^ data_out[275] ^ data_out[274] ^ data_out[273] ^ data_out[272] ^ data_out[271] ^ data_out[270] ^ data_out[269] ^ data_out[268] ^ data_out[267] ^ data_out[266] ^ data_out[265] ^ data_out[264] ^ data_out[263] ^ data_out[262] ^ data_out[261] ^ data_out[260] ^ data_out[259] ^ data_out[258] ^ data_out[257] ^ data_out[256] ^ data_out[255] ^ data_out[127] ^ data_out[126] ^ data_out[125] ^ data_out[124] ^ data_out[123] ^ data_out[122] ^ data_out[121] ^ data_out[120] ^ data_out[119] ^ data_out[118] ^ data_out[117] ^ data_out[116] ^ data_out[115] ^ data_out[114] ^ data_out[113] ^ data_out[112] ^ data_out[111] ^ data_out[110] ^ data_out[109] ^ data_out[108] ^ data_out[107] ^ data_out[106] ^ data_out[105] ^ data_out[104] ^ data_out[103] ^ data_out[102] ^ data_out[101] ^ data_out[100] ^ data_out[99] ^ data_out[98] ^ data_out[97] ^ data_out[96] ^ data_out[95] ^ data_out[94] ^ data_out[93] ^ data_out[92] ^ data_out[91] ^ data_out[90] ^ data_out[89] ^ data_out[88] ^ data_out[87] ^ data_out[86] ^ data_out[85] ^ data_out[84] ^ data_out[83] ^ data_out[82] ^ data_out[81] ^ data_out[80] ^ data_out[79] ^ data_out[78] ^ data_out[77] ^ data_out[76] ^ data_out[75] ^ data_out[74] ^ data_out[73] ^ data_out[72] ^ data_out[71] ^ data_out[70] ^ data_out[69] ^ data_out[68] ^ data_out[67] ^ data_out[66] ^ data_out[65] ^ data_out[64] ^ data_out[63] ^ data_out[62] ^ data_out[61] ^ data_out[60] ^ data_out[59] ^ data_out[58] ^ data_out[57] ^ data_out[56] ^ data_out[55] ^ data_out[54] ^ data_out[53] ^ data_out[52] ^ data_out[51] ^ data_out[50] ^ data_out[49] ^ data_out[48] ^ data_out[47] ^ data_out[46] ^ data_out[45] ^ data_out[44] ^ data_out[43] ^ data_out[42] ^ data_out[41] ^ data_out[40] ^ data_out[39] ^ data_out[38] ^ data_out[37] ^ data_out[36] ^ data_out[35] ^ data_out[34] ^ data_out[33] ^ data_out[32] ^ data_out[31] ^ data_out[30] ^ data_out[29] ^ data_out[28] ^ data_out[27] ^ data_out[26] ^ data_out[25] ^ data_out[24] ^ data_out[23] ^ data_out[22] ^ data_out[21] ^ data_out[20] ^ data_out[19] ^ data_out[18] ^ data_out[17] ^ data_out[16] ^ data_out[15] ^ data_out[14] ^ data_out[13] ^ data_out[12] ^ data_out[11] ^ data_out[10] ^ data_out[9] ^ data_out[8] ^ data_out[7] ^ data_out[6] ^ data_out[5] ^ data_out[4] ^ data_out[3] ^ data_out[2] ^ data_out[1] ^ data_out[0] ^ checker_out[7] ;
    syndrome[8] = data_out[254] ^ data_out[253] ^ data_out[252] ^ data_out[251] ^ data_out[250] ^ data_out[249] ^ data_out[248] ^ data_out[247] ^ data_out[246] ^ data_out[245] ^ data_out[244] ^ data_out[243] ^ data_out[242] ^ data_out[241] ^ data_out[240] ^ data_out[239] ^ data_out[238] ^ data_out[237] ^ data_out[236] ^ data_out[235] ^ data_out[234] ^ data_out[233] ^ data_out[232] ^ data_out[231] ^ data_out[230] ^ data_out[229] ^ data_out[228] ^ data_out[227] ^ data_out[226] ^ data_out[225] ^ data_out[224] ^ data_out[223] ^ data_out[222] ^ data_out[221] ^ data_out[220] ^ data_out[219] ^ data_out[218] ^ data_out[217] ^ data_out[216] ^ data_out[215] ^ data_out[214] ^ data_out[213] ^ data_out[212] ^ data_out[211] ^ data_out[210] ^ data_out[209] ^ data_out[208] ^ data_out[207] ^ data_out[206] ^ data_out[205] ^ data_out[204] ^ data_out[203] ^ data_out[202] ^ data_out[201] ^ data_out[200] ^ data_out[199] ^ data_out[198] ^ data_out[197] ^ data_out[196] ^ data_out[195] ^ data_out[194] ^ data_out[193] ^ data_out[192] ^ data_out[191] ^ data_out[190] ^ data_out[189] ^ data_out[188] ^ data_out[187] ^ data_out[186] ^ data_out[185] ^ data_out[184] ^ data_out[183] ^ data_out[182] ^ data_out[181] ^ data_out[180] ^ data_out[179] ^ data_out[178] ^ data_out[177] ^ data_out[176] ^ data_out[175] ^ data_out[174] ^ data_out[173] ^ data_out[172] ^ data_out[171] ^ data_out[170] ^ data_out[169] ^ data_out[168] ^ data_out[167] ^ data_out[166] ^ data_out[165] ^ data_out[164] ^ data_out[163] ^ data_out[162] ^ data_out[161] ^ data_out[160] ^ data_out[159] ^ data_out[158] ^ data_out[157] ^ data_out[156] ^ data_out[155] ^ data_out[154] ^ data_out[153] ^ data_out[152] ^ data_out[151] ^ data_out[150] ^ data_out[149] ^ data_out[148] ^ data_out[147] ^ data_out[146] ^ data_out[145] ^ data_out[144] ^ data_out[143] ^ data_out[142] ^ data_out[141] ^ data_out[140] ^ data_out[139] ^ data_out[138] ^ data_out[137] ^ data_out[136] ^ data_out[135] ^ data_out[134] ^ data_out[133] ^ data_out[132] ^ data_out[131] ^ data_out[130] ^ data_out[129] ^ data_out[128] ^ data_out[127] ^ data_out[126] ^ data_out[125] ^ data_out[124] ^ data_out[123] ^ data_out[122] ^ data_out[121] ^ data_out[120] ^ data_out[119] ^ data_out[118] ^ data_out[117] ^ data_out[116] ^ data_out[115] ^ data_out[114] ^ data_out[113] ^ data_out[112] ^ data_out[111] ^ data_out[110] ^ data_out[109] ^ data_out[108] ^ data_out[107] ^ data_out[106] ^ data_out[105] ^ data_out[104] ^ data_out[103] ^ data_out[102] ^ data_out[101] ^ data_out[100] ^ data_out[99] ^ data_out[98] ^ data_out[97] ^ data_out[96] ^ data_out[95] ^ data_out[94] ^ data_out[93] ^ data_out[92] ^ data_out[91] ^ data_out[90] ^ data_out[89] ^ data_out[88] ^ data_out[87] ^ data_out[86] ^ data_out[85] ^ data_out[84] ^ data_out[83] ^ data_out[82] ^ data_out[81] ^ data_out[80] ^ data_out[79] ^ data_out[78] ^ data_out[77] ^ data_out[76] ^ data_out[75] ^ data_out[74] ^ data_out[73] ^ data_out[72] ^ data_out[71] ^ data_out[70] ^ data_out[69] ^ data_out[68] ^ data_out[67] ^ data_out[66] ^ data_out[65] ^ data_out[64] ^ data_out[63] ^ data_out[62] ^ data_out[61] ^ data_out[60] ^ data_out[59] ^ data_out[58] ^ data_out[57] ^ data_out[56] ^ data_out[55] ^ data_out[54] ^ data_out[53] ^ data_out[52] ^ data_out[51] ^ data_out[50] ^ data_out[49] ^ data_out[48] ^ data_out[47] ^ data_out[46] ^ data_out[45] ^ data_out[44] ^ data_out[43] ^ data_out[42] ^ data_out[41] ^ data_out[40] ^ data_out[39] ^ data_out[38] ^ data_out[37] ^ data_out[36] ^ data_out[35] ^ data_out[34] ^ data_out[33] ^ data_out[32] ^ data_out[31] ^ data_out[30] ^ data_out[29] ^ data_out[28] ^ data_out[27] ^ data_out[26] ^ data_out[25] ^ data_out[24] ^ data_out[23] ^ data_out[22] ^ data_out[21] ^ data_out[20] ^ data_out[19] ^ data_out[18] ^ data_out[17] ^ data_out[16] ^ data_out[15] ^ data_out[14] ^ data_out[13] ^ data_out[12] ^ data_out[11] ^ data_out[10] ^ data_out[9] ^ data_out[8] ^ data_out[7] ^ data_out[6] ^ data_out[5] ^ data_out[4] ^ data_out[3] ^ data_out[2] ^ data_out[1] ^ data_out[0] ^ checker_out[8] ;

    parity = data_out[0] ^ data_out[1] ^ data_out[2] ^ data_out[3] ^ data_out[4] ^ data_out[5] ^ data_out[6] ^ data_out[7] ^ data_out[8] ^ data_out[9] ^ data_out[10] ^ data_out[11] ^ data_out[12] ^ data_out[13] ^ data_out[14] ^ data_out[15] ^ data_out[16] ^ data_out[17] ^ data_out[18] ^ data_out[19] ^ data_out[20] ^ data_out[21] ^ data_out[22] ^ data_out[23] ^ data_out[24] ^ data_out[25] ^ data_out[26] ^ data_out[27] ^ data_out[28] ^ data_out[29] ^ data_out[30] ^ data_out[31] ^ data_out[32] ^ data_out[33] ^ data_out[34] ^ data_out[35] ^ data_out[36] ^ data_out[37] ^ data_out[38] ^ data_out[39] ^ data_out[40] ^ data_out[41] ^ data_out[42] ^ data_out[43] ^ data_out[44] ^ data_out[45] ^ data_out[46] ^ data_out[47] ^ data_out[48] ^ data_out[49] ^ data_out[50] ^ data_out[51] ^ data_out[52] ^ data_out[53] ^ data_out[54] ^ data_out[55] ^ data_out[56] ^ data_out[57] ^ data_out[58] ^ data_out[59] ^ data_out[60] ^ data_out[61] ^ data_out[62] ^ data_out[63] ^ data_out[64] ^ data_out[65] ^ data_out[66] ^ data_out[67] ^ data_out[68] ^ data_out[69] ^ data_out[70] ^ data_out[71] ^ data_out[72] ^ data_out[73] ^ data_out[74] ^ data_out[75] ^ data_out[76] ^ data_out[77] ^ data_out[78] ^ data_out[79] ^ data_out[80] ^ data_out[81] ^ data_out[82] ^ data_out[83] ^ data_out[84] ^ data_out[85] ^ data_out[86] ^ data_out[87] ^ data_out[88] ^ data_out[89] ^ data_out[90] ^ data_out[91] ^ data_out[92] ^ data_out[93] ^ data_out[94] ^ data_out[95] ^ data_out[96] ^ data_out[97] ^ data_out[98] ^ data_out[99] ^ data_out[100] ^ data_out[101] ^ data_out[102] ^ data_out[103] ^ data_out[104] ^ data_out[105] ^ data_out[106] ^ data_out[107] ^ data_out[108] ^ data_out[109] ^ data_out[110] ^ data_out[111] ^ data_out[112] ^ data_out[113] ^ data_out[114] ^ data_out[115] ^ data_out[116] ^ data_out[117] ^ data_out[118] ^ data_out[119] ^ data_out[120] ^ data_out[121] ^ data_out[122] ^ data_out[123] ^ data_out[124] ^ data_out[125] ^ data_out[126] ^ data_out[127] ^ data_out[128] ^ data_out[129] ^ data_out[130] ^ data_out[131] ^ data_out[132] ^ data_out[133] ^ data_out[134] ^ data_out[135] ^ data_out[136] ^ data_out[137] ^ data_out[138] ^ data_out[139] ^ data_out[140] ^ data_out[141] ^ data_out[142] ^ data_out[143] ^ data_out[144] ^ data_out[145] ^ data_out[146] ^ data_out[147] ^ data_out[148] ^ data_out[149] ^ data_out[150] ^ data_out[151] ^ data_out[152] ^ data_out[153] ^ data_out[154] ^ data_out[155] ^ data_out[156] ^ data_out[157] ^ data_out[158] ^ data_out[159] ^ data_out[160] ^ data_out[161] ^ data_out[162] ^ data_out[163] ^ data_out[164] ^ data_out[165] ^ data_out[166] ^ data_out[167] ^ data_out[168] ^ data_out[169] ^ data_out[170] ^ data_out[171] ^ data_out[172] ^ data_out[173] ^ data_out[174] ^ data_out[175] ^ data_out[176] ^ data_out[177] ^ data_out[178] ^ data_out[179] ^ data_out[180] ^ data_out[181] ^ data_out[182] ^ data_out[183] ^ data_out[184] ^ data_out[185] ^ data_out[186] ^ data_out[187] ^ data_out[188] ^ data_out[189] ^ data_out[190] ^ data_out[191] ^ data_out[192] ^ data_out[193] ^ data_out[194] ^ data_out[195] ^ data_out[196] ^ data_out[197] ^ data_out[198] ^ data_out[199] ^ data_out[200] ^ data_out[201] ^ data_out[202] ^ data_out[203] ^ data_out[204] ^ data_out[205] ^ data_out[206] ^ data_out[207] ^ data_out[208] ^ data_out[209] ^ data_out[210] ^ data_out[211] ^ data_out[212] ^ data_out[213] ^ data_out[214] ^ data_out[215] ^ data_out[216] ^ data_out[217] ^ data_out[218] ^ data_out[219] ^ data_out[220] ^ data_out[221] ^ data_out[222] ^ data_out[223] ^ data_out[224] ^ data_out[225] ^ data_out[226] ^ data_out[227] ^ data_out[228] ^ data_out[229] ^ data_out[230] ^ data_out[231] ^ data_out[232] ^ data_out[233] ^ data_out[234] ^ data_out[235] ^ data_out[236] ^ data_out[237] ^ data_out[238] ^ data_out[239] ^ data_out[240] ^ data_out[241] ^ data_out[242] ^ data_out[243] ^ data_out[244] ^ data_out[245] ^ data_out[246] ^ data_out[247] ^ data_out[248] ^ data_out[249] ^ data_out[250] ^ data_out[251] ^ data_out[252] ^ data_out[253] ^ data_out[254] ^ data_out[255] ^ data_out[256] ^ data_out[257] ^ data_out[258] ^ data_out[259] ^ data_out[260] ^ data_out[261] ^ data_out[262] ^ data_out[263] ^ data_out[264] ^ data_out[265] ^ data_out[266] ^ data_out[267] ^ data_out[268] ^ data_out[269] ^ data_out[270] ^ data_out[271] ^ data_out[272] ^ data_out[273] ^ data_out[274] ^ data_out[275] ^ data_out[276] ^ data_out[277] ^ data_out[278] ^ data_out[279] ^ data_out[280] ^ data_out[281] ^ data_out[282] ^ data_out[283] ^ data_out[284] ^ data_out[285] ^ data_out[286] ^ data_out[287] ^ data_out[288] ^ data_out[289] ^ data_out[290] ^ data_out[291] ^ data_out[292] ^ data_out[293] ^ data_out[294] ^ data_out[295] ^ data_out[296] ^ data_out[297] ^ data_out[298] ^ data_out[299] ^ data_out[300] ^ data_out[301] ^ data_out[302] ^ data_out[303] ^ data_out[304] ^ data_out[305] ^ data_out[306] ^ data_out[307] ^ data_out[308] ^ data_out[309] ^ data_out[310] ^ data_out[311] ^ data_out[312] ^ data_out[313] ^ data_out[314] ^ data_out[315] ^ data_out[316] ^ data_out[317] ^ data_out[318] ^ data_out[319] ^ data_out[320] ^ data_out[321] ^ data_out[322] ^ data_out[323] ^ data_out[324] ^ data_out[325] ^ data_out[326] ^ data_out[327] ^ data_out[328] ^ data_out[329] ^ data_out[330] ^ data_out[331] ^ data_out[332] ^ data_out[333] ^ data_out[334] ^ data_out[335] ^ data_out[336] ^ data_out[337] ^ data_out[338] ^ data_out[339] ^ data_out[340] ^ data_out[341] ^ data_out[342] ^ data_out[343] ^ data_out[344] ^ data_out[345] ^ data_out[346] ^ data_out[347] ^ data_out[348] ^ data_out[349] ^ data_out[350] ^ data_out[351] ^ data_out[352] ^ data_out[353] ^ data_out[354] ^ data_out[355] ^ data_out[356] ^ data_out[357] ^ data_out[358] ^ data_out[359] ^ data_out[360] ^ data_out[361] ^ data_out[362] ^ data_out[363] ^ data_out[364] ^ data_out[365] ^ data_out[366] ^ data_out[367] ^ data_out[368] ^ data_out[369] ^ data_out[370] ^ data_out[371] ^ data_out[372] ^ data_out[373] ^ data_out[374] ^ data_out[375] ^ data_out[376] ^ data_out[377] ^ data_out[378] ^ data_out[379] ^ data_out[380] ^ data_out[381] ^ data_out[382] ^ data_out[383] ^ data_out[384] ^ data_out[385] ^ data_out[386] ^ data_out[387] ^ data_out[388] ^ data_out[389] ^ data_out[390] ^ data_out[391] ^ data_out[392] ^ data_out[393] ^ data_out[394] ^ data_out[395] ^ data_out[396] ^ data_out[397] ^ data_out[398] ^ data_out[399] ^ data_out[400] ^ data_out[401] ^ data_out[402] ^ data_out[403] ^ data_out[404] ^ data_out[405] ^ data_out[406] ^ data_out[407] ^ data_out[408] ^ data_out[409] ^ data_out[410] ^ data_out[411] ^ data_out[412] ^ data_out[413] ^ data_out[414] ^ data_out[415] ^ data_out[416] ^ data_out[417] ^ data_out[418] ^ data_out[419] ^ data_out[420] ^ data_out[421] ^ data_out[422] ^ data_out[423] ^ data_out[424] ^ data_out[425] ^ data_out[426] ^ data_out[427] ^ data_out[428] ^ data_out[429] ^ data_out[430] ^ data_out[431] ^ data_out[432] ^ data_out[433] ^ data_out[434] ^ data_out[435] ^ data_out[436] ^ data_out[437] ^ data_out[438] ^ data_out[439] ^ data_out[440] ^ data_out[441] ^ data_out[442] ^ data_out[443] ^ data_out[444] ^ data_out[445] ^ data_out[446] ^ data_out[447] ^ data_out[448] ^ data_out[449] ^ data_out[450] ^ data_out[451] ^ data_out[452] ^ data_out[453] ^ data_out[454] ^ data_out[455] ^ data_out[456] ^ data_out[457] ^ data_out[458] ^ data_out[459] ^ data_out[460] ^ data_out[461] ^ data_out[462] ^ data_out[463] ^ data_out[464] ^ data_out[465] ^ data_out[466] ^ data_out[467] ^ data_out[468] ^ data_out[469] ^ data_out[470] ^ data_out[471] ^ data_out[472] ^ data_out[473] ^ data_out[474] ^ data_out[475] ^ data_out[476] ^ data_out[477] ^ data_out[478] ^ data_out[479] ^ data_out[480] ^ data_out[481] ^ data_out[482] ^ data_out[483] ^ data_out[484] ^ data_out[485] ^ data_out[486] ^ data_out[487] ^ data_out[488] ^ data_out[489] ^ data_out[490] ^ data_out[491] ^ data_out[492] ^ data_out[493] ^ data_out[494] ^ data_out[495] ^ data_out[496] ^ data_out[497] ^ data_out[498] ^ data_out[499] ^ data_out[500] ^ data_out[501] ^ checker_out[0] ^ checker_out[1] ^ checker_out[2] ^ checker_out[3] ^ checker_out[4] ^ checker_out[5] ^ checker_out[6] ^ checker_out[7] ^ checker_out[8] ^ parity_out ;

    error = 0;
    if (syndrome == 0 && parity == 0) begin
        error = 0;
    end
    if (syndrome != 0 && parity == 0) begin
        error = 1;
    end
    if (syndrome == 0 && parity != 0) begin
        error = 0;
    end
    if (syndrome != 0 && parity != 0) begin
        error = 0;
    end

    correct_data_out = data_out;
    if (error == 0 && syndrome != 0) begin
        case(syndrome)
            3: correct_data_out[501] = ~data_out[501];
            5: correct_data_out[500] = ~data_out[500];
            6: correct_data_out[499] = ~data_out[499];
            7: correct_data_out[498] = ~data_out[498];
            9: correct_data_out[497] = ~data_out[497];
            10: correct_data_out[496] = ~data_out[496];
            11: correct_data_out[495] = ~data_out[495];
            12: correct_data_out[494] = ~data_out[494];
            13: correct_data_out[493] = ~data_out[493];
            14: correct_data_out[492] = ~data_out[492];
            15: correct_data_out[491] = ~data_out[491];
            17: correct_data_out[490] = ~data_out[490];
            18: correct_data_out[489] = ~data_out[489];
            19: correct_data_out[488] = ~data_out[488];
            20: correct_data_out[487] = ~data_out[487];
            21: correct_data_out[486] = ~data_out[486];
            22: correct_data_out[485] = ~data_out[485];
            23: correct_data_out[484] = ~data_out[484];
            24: correct_data_out[483] = ~data_out[483];
            25: correct_data_out[482] = ~data_out[482];
            26: correct_data_out[481] = ~data_out[481];
            27: correct_data_out[480] = ~data_out[480];
            28: correct_data_out[479] = ~data_out[479];
            29: correct_data_out[478] = ~data_out[478];
            30: correct_data_out[477] = ~data_out[477];
            31: correct_data_out[476] = ~data_out[476];
            33: correct_data_out[475] = ~data_out[475];
            34: correct_data_out[474] = ~data_out[474];
            35: correct_data_out[473] = ~data_out[473];
            36: correct_data_out[472] = ~data_out[472];
            37: correct_data_out[471] = ~data_out[471];
            38: correct_data_out[470] = ~data_out[470];
            39: correct_data_out[469] = ~data_out[469];
            40: correct_data_out[468] = ~data_out[468];
            41: correct_data_out[467] = ~data_out[467];
            42: correct_data_out[466] = ~data_out[466];
            43: correct_data_out[465] = ~data_out[465];
            44: correct_data_out[464] = ~data_out[464];
            45: correct_data_out[463] = ~data_out[463];
            46: correct_data_out[462] = ~data_out[462];
            47: correct_data_out[461] = ~data_out[461];
            48: correct_data_out[460] = ~data_out[460];
            49: correct_data_out[459] = ~data_out[459];
            50: correct_data_out[458] = ~data_out[458];
            51: correct_data_out[457] = ~data_out[457];
            52: correct_data_out[456] = ~data_out[456];
            53: correct_data_out[455] = ~data_out[455];
            54: correct_data_out[454] = ~data_out[454];
            55: correct_data_out[453] = ~data_out[453];
            56: correct_data_out[452] = ~data_out[452];
            57: correct_data_out[451] = ~data_out[451];
            58: correct_data_out[450] = ~data_out[450];
            59: correct_data_out[449] = ~data_out[449];
            60: correct_data_out[448] = ~data_out[448];
            61: correct_data_out[447] = ~data_out[447];
            62: correct_data_out[446] = ~data_out[446];
            63: correct_data_out[445] = ~data_out[445];
            65: correct_data_out[444] = ~data_out[444];
            66: correct_data_out[443] = ~data_out[443];
            67: correct_data_out[442] = ~data_out[442];
            68: correct_data_out[441] = ~data_out[441];
            69: correct_data_out[440] = ~data_out[440];
            70: correct_data_out[439] = ~data_out[439];
            71: correct_data_out[438] = ~data_out[438];
            72: correct_data_out[437] = ~data_out[437];
            73: correct_data_out[436] = ~data_out[436];
            74: correct_data_out[435] = ~data_out[435];
            75: correct_data_out[434] = ~data_out[434];
            76: correct_data_out[433] = ~data_out[433];
            77: correct_data_out[432] = ~data_out[432];
            78: correct_data_out[431] = ~data_out[431];
            79: correct_data_out[430] = ~data_out[430];
            80: correct_data_out[429] = ~data_out[429];
            81: correct_data_out[428] = ~data_out[428];
            82: correct_data_out[427] = ~data_out[427];
            83: correct_data_out[426] = ~data_out[426];
            84: correct_data_out[425] = ~data_out[425];
            85: correct_data_out[424] = ~data_out[424];
            86: correct_data_out[423] = ~data_out[423];
            87: correct_data_out[422] = ~data_out[422];
            88: correct_data_out[421] = ~data_out[421];
            89: correct_data_out[420] = ~data_out[420];
            90: correct_data_out[419] = ~data_out[419];
            91: correct_data_out[418] = ~data_out[418];
            92: correct_data_out[417] = ~data_out[417];
            93: correct_data_out[416] = ~data_out[416];
            94: correct_data_out[415] = ~data_out[415];
            95: correct_data_out[414] = ~data_out[414];
            96: correct_data_out[413] = ~data_out[413];
            97: correct_data_out[412] = ~data_out[412];
            98: correct_data_out[411] = ~data_out[411];
            99: correct_data_out[410] = ~data_out[410];
            100: correct_data_out[409] = ~data_out[409];
            101: correct_data_out[408] = ~data_out[408];
            102: correct_data_out[407] = ~data_out[407];
            103: correct_data_out[406] = ~data_out[406];
            104: correct_data_out[405] = ~data_out[405];
            105: correct_data_out[404] = ~data_out[404];
            106: correct_data_out[403] = ~data_out[403];
            107: correct_data_out[402] = ~data_out[402];
            108: correct_data_out[401] = ~data_out[401];
            109: correct_data_out[400] = ~data_out[400];
            110: correct_data_out[399] = ~data_out[399];
            111: correct_data_out[398] = ~data_out[398];
            112: correct_data_out[397] = ~data_out[397];
            113: correct_data_out[396] = ~data_out[396];
            114: correct_data_out[395] = ~data_out[395];
            115: correct_data_out[394] = ~data_out[394];
            116: correct_data_out[393] = ~data_out[393];
            117: correct_data_out[392] = ~data_out[392];
            118: correct_data_out[391] = ~data_out[391];
            119: correct_data_out[390] = ~data_out[390];
            120: correct_data_out[389] = ~data_out[389];
            121: correct_data_out[388] = ~data_out[388];
            122: correct_data_out[387] = ~data_out[387];
            123: correct_data_out[386] = ~data_out[386];
            124: correct_data_out[385] = ~data_out[385];
            125: correct_data_out[384] = ~data_out[384];
            126: correct_data_out[383] = ~data_out[383];
            127: correct_data_out[382] = ~data_out[382];
            129: correct_data_out[381] = ~data_out[381];
            130: correct_data_out[380] = ~data_out[380];
            131: correct_data_out[379] = ~data_out[379];
            132: correct_data_out[378] = ~data_out[378];
            133: correct_data_out[377] = ~data_out[377];
            134: correct_data_out[376] = ~data_out[376];
            135: correct_data_out[375] = ~data_out[375];
            136: correct_data_out[374] = ~data_out[374];
            137: correct_data_out[373] = ~data_out[373];
            138: correct_data_out[372] = ~data_out[372];
            139: correct_data_out[371] = ~data_out[371];
            140: correct_data_out[370] = ~data_out[370];
            141: correct_data_out[369] = ~data_out[369];
            142: correct_data_out[368] = ~data_out[368];
            143: correct_data_out[367] = ~data_out[367];
            144: correct_data_out[366] = ~data_out[366];
            145: correct_data_out[365] = ~data_out[365];
            146: correct_data_out[364] = ~data_out[364];
            147: correct_data_out[363] = ~data_out[363];
            148: correct_data_out[362] = ~data_out[362];
            149: correct_data_out[361] = ~data_out[361];
            150: correct_data_out[360] = ~data_out[360];
            151: correct_data_out[359] = ~data_out[359];
            152: correct_data_out[358] = ~data_out[358];
            153: correct_data_out[357] = ~data_out[357];
            154: correct_data_out[356] = ~data_out[356];
            155: correct_data_out[355] = ~data_out[355];
            156: correct_data_out[354] = ~data_out[354];
            157: correct_data_out[353] = ~data_out[353];
            158: correct_data_out[352] = ~data_out[352];
            159: correct_data_out[351] = ~data_out[351];
            160: correct_data_out[350] = ~data_out[350];
            161: correct_data_out[349] = ~data_out[349];
            162: correct_data_out[348] = ~data_out[348];
            163: correct_data_out[347] = ~data_out[347];
            164: correct_data_out[346] = ~data_out[346];
            165: correct_data_out[345] = ~data_out[345];
            166: correct_data_out[344] = ~data_out[344];
            167: correct_data_out[343] = ~data_out[343];
            168: correct_data_out[342] = ~data_out[342];
            169: correct_data_out[341] = ~data_out[341];
            170: correct_data_out[340] = ~data_out[340];
            171: correct_data_out[339] = ~data_out[339];
            172: correct_data_out[338] = ~data_out[338];
            173: correct_data_out[337] = ~data_out[337];
            174: correct_data_out[336] = ~data_out[336];
            175: correct_data_out[335] = ~data_out[335];
            176: correct_data_out[334] = ~data_out[334];
            177: correct_data_out[333] = ~data_out[333];
            178: correct_data_out[332] = ~data_out[332];
            179: correct_data_out[331] = ~data_out[331];
            180: correct_data_out[330] = ~data_out[330];
            181: correct_data_out[329] = ~data_out[329];
            182: correct_data_out[328] = ~data_out[328];
            183: correct_data_out[327] = ~data_out[327];
            184: correct_data_out[326] = ~data_out[326];
            185: correct_data_out[325] = ~data_out[325];
            186: correct_data_out[324] = ~data_out[324];
            187: correct_data_out[323] = ~data_out[323];
            188: correct_data_out[322] = ~data_out[322];
            189: correct_data_out[321] = ~data_out[321];
            190: correct_data_out[320] = ~data_out[320];
            191: correct_data_out[319] = ~data_out[319];
            192: correct_data_out[318] = ~data_out[318];
            193: correct_data_out[317] = ~data_out[317];
            194: correct_data_out[316] = ~data_out[316];
            195: correct_data_out[315] = ~data_out[315];
            196: correct_data_out[314] = ~data_out[314];
            197: correct_data_out[313] = ~data_out[313];
            198: correct_data_out[312] = ~data_out[312];
            199: correct_data_out[311] = ~data_out[311];
            200: correct_data_out[310] = ~data_out[310];
            201: correct_data_out[309] = ~data_out[309];
            202: correct_data_out[308] = ~data_out[308];
            203: correct_data_out[307] = ~data_out[307];
            204: correct_data_out[306] = ~data_out[306];
            205: correct_data_out[305] = ~data_out[305];
            206: correct_data_out[304] = ~data_out[304];
            207: correct_data_out[303] = ~data_out[303];
            208: correct_data_out[302] = ~data_out[302];
            209: correct_data_out[301] = ~data_out[301];
            210: correct_data_out[300] = ~data_out[300];
            211: correct_data_out[299] = ~data_out[299];
            212: correct_data_out[298] = ~data_out[298];
            213: correct_data_out[297] = ~data_out[297];
            214: correct_data_out[296] = ~data_out[296];
            215: correct_data_out[295] = ~data_out[295];
            216: correct_data_out[294] = ~data_out[294];
            217: correct_data_out[293] = ~data_out[293];
            218: correct_data_out[292] = ~data_out[292];
            219: correct_data_out[291] = ~data_out[291];
            220: correct_data_out[290] = ~data_out[290];
            221: correct_data_out[289] = ~data_out[289];
            222: correct_data_out[288] = ~data_out[288];
            223: correct_data_out[287] = ~data_out[287];
            224: correct_data_out[286] = ~data_out[286];
            225: correct_data_out[285] = ~data_out[285];
            226: correct_data_out[284] = ~data_out[284];
            227: correct_data_out[283] = ~data_out[283];
            228: correct_data_out[282] = ~data_out[282];
            229: correct_data_out[281] = ~data_out[281];
            230: correct_data_out[280] = ~data_out[280];
            231: correct_data_out[279] = ~data_out[279];
            232: correct_data_out[278] = ~data_out[278];
            233: correct_data_out[277] = ~data_out[277];
            234: correct_data_out[276] = ~data_out[276];
            235: correct_data_out[275] = ~data_out[275];
            236: correct_data_out[274] = ~data_out[274];
            237: correct_data_out[273] = ~data_out[273];
            238: correct_data_out[272] = ~data_out[272];
            239: correct_data_out[271] = ~data_out[271];
            240: correct_data_out[270] = ~data_out[270];
            241: correct_data_out[269] = ~data_out[269];
            242: correct_data_out[268] = ~data_out[268];
            243: correct_data_out[267] = ~data_out[267];
            244: correct_data_out[266] = ~data_out[266];
            245: correct_data_out[265] = ~data_out[265];
            246: correct_data_out[264] = ~data_out[264];
            247: correct_data_out[263] = ~data_out[263];
            248: correct_data_out[262] = ~data_out[262];
            249: correct_data_out[261] = ~data_out[261];
            250: correct_data_out[260] = ~data_out[260];
            251: correct_data_out[259] = ~data_out[259];
            252: correct_data_out[258] = ~data_out[258];
            253: correct_data_out[257] = ~data_out[257];
            254: correct_data_out[256] = ~data_out[256];
            255: correct_data_out[255] = ~data_out[255];
            257: correct_data_out[254] = ~data_out[254];
            258: correct_data_out[253] = ~data_out[253];
            259: correct_data_out[252] = ~data_out[252];
            260: correct_data_out[251] = ~data_out[251];
            261: correct_data_out[250] = ~data_out[250];
            262: correct_data_out[249] = ~data_out[249];
            263: correct_data_out[248] = ~data_out[248];
            264: correct_data_out[247] = ~data_out[247];
            265: correct_data_out[246] = ~data_out[246];
            266: correct_data_out[245] = ~data_out[245];
            267: correct_data_out[244] = ~data_out[244];
            268: correct_data_out[243] = ~data_out[243];
            269: correct_data_out[242] = ~data_out[242];
            270: correct_data_out[241] = ~data_out[241];
            271: correct_data_out[240] = ~data_out[240];
            272: correct_data_out[239] = ~data_out[239];
            273: correct_data_out[238] = ~data_out[238];
            274: correct_data_out[237] = ~data_out[237];
            275: correct_data_out[236] = ~data_out[236];
            276: correct_data_out[235] = ~data_out[235];
            277: correct_data_out[234] = ~data_out[234];
            278: correct_data_out[233] = ~data_out[233];
            279: correct_data_out[232] = ~data_out[232];
            280: correct_data_out[231] = ~data_out[231];
            281: correct_data_out[230] = ~data_out[230];
            282: correct_data_out[229] = ~data_out[229];
            283: correct_data_out[228] = ~data_out[228];
            284: correct_data_out[227] = ~data_out[227];
            285: correct_data_out[226] = ~data_out[226];
            286: correct_data_out[225] = ~data_out[225];
            287: correct_data_out[224] = ~data_out[224];
            288: correct_data_out[223] = ~data_out[223];
            289: correct_data_out[222] = ~data_out[222];
            290: correct_data_out[221] = ~data_out[221];
            291: correct_data_out[220] = ~data_out[220];
            292: correct_data_out[219] = ~data_out[219];
            293: correct_data_out[218] = ~data_out[218];
            294: correct_data_out[217] = ~data_out[217];
            295: correct_data_out[216] = ~data_out[216];
            296: correct_data_out[215] = ~data_out[215];
            297: correct_data_out[214] = ~data_out[214];
            298: correct_data_out[213] = ~data_out[213];
            299: correct_data_out[212] = ~data_out[212];
            300: correct_data_out[211] = ~data_out[211];
            301: correct_data_out[210] = ~data_out[210];
            302: correct_data_out[209] = ~data_out[209];
            303: correct_data_out[208] = ~data_out[208];
            304: correct_data_out[207] = ~data_out[207];
            305: correct_data_out[206] = ~data_out[206];
            306: correct_data_out[205] = ~data_out[205];
            307: correct_data_out[204] = ~data_out[204];
            308: correct_data_out[203] = ~data_out[203];
            309: correct_data_out[202] = ~data_out[202];
            310: correct_data_out[201] = ~data_out[201];
            311: correct_data_out[200] = ~data_out[200];
            312: correct_data_out[199] = ~data_out[199];
            313: correct_data_out[198] = ~data_out[198];
            314: correct_data_out[197] = ~data_out[197];
            315: correct_data_out[196] = ~data_out[196];
            316: correct_data_out[195] = ~data_out[195];
            317: correct_data_out[194] = ~data_out[194];
            318: correct_data_out[193] = ~data_out[193];
            319: correct_data_out[192] = ~data_out[192];
            320: correct_data_out[191] = ~data_out[191];
            321: correct_data_out[190] = ~data_out[190];
            322: correct_data_out[189] = ~data_out[189];
            323: correct_data_out[188] = ~data_out[188];
            324: correct_data_out[187] = ~data_out[187];
            325: correct_data_out[186] = ~data_out[186];
            326: correct_data_out[185] = ~data_out[185];
            327: correct_data_out[184] = ~data_out[184];
            328: correct_data_out[183] = ~data_out[183];
            329: correct_data_out[182] = ~data_out[182];
            330: correct_data_out[181] = ~data_out[181];
            331: correct_data_out[180] = ~data_out[180];
            332: correct_data_out[179] = ~data_out[179];
            333: correct_data_out[178] = ~data_out[178];
            334: correct_data_out[177] = ~data_out[177];
            335: correct_data_out[176] = ~data_out[176];
            336: correct_data_out[175] = ~data_out[175];
            337: correct_data_out[174] = ~data_out[174];
            338: correct_data_out[173] = ~data_out[173];
            339: correct_data_out[172] = ~data_out[172];
            340: correct_data_out[171] = ~data_out[171];
            341: correct_data_out[170] = ~data_out[170];
            342: correct_data_out[169] = ~data_out[169];
            343: correct_data_out[168] = ~data_out[168];
            344: correct_data_out[167] = ~data_out[167];
            345: correct_data_out[166] = ~data_out[166];
            346: correct_data_out[165] = ~data_out[165];
            347: correct_data_out[164] = ~data_out[164];
            348: correct_data_out[163] = ~data_out[163];
            349: correct_data_out[162] = ~data_out[162];
            350: correct_data_out[161] = ~data_out[161];
            351: correct_data_out[160] = ~data_out[160];
            352: correct_data_out[159] = ~data_out[159];
            353: correct_data_out[158] = ~data_out[158];
            354: correct_data_out[157] = ~data_out[157];
            355: correct_data_out[156] = ~data_out[156];
            356: correct_data_out[155] = ~data_out[155];
            357: correct_data_out[154] = ~data_out[154];
            358: correct_data_out[153] = ~data_out[153];
            359: correct_data_out[152] = ~data_out[152];
            360: correct_data_out[151] = ~data_out[151];
            361: correct_data_out[150] = ~data_out[150];
            362: correct_data_out[149] = ~data_out[149];
            363: correct_data_out[148] = ~data_out[148];
            364: correct_data_out[147] = ~data_out[147];
            365: correct_data_out[146] = ~data_out[146];
            366: correct_data_out[145] = ~data_out[145];
            367: correct_data_out[144] = ~data_out[144];
            368: correct_data_out[143] = ~data_out[143];
            369: correct_data_out[142] = ~data_out[142];
            370: correct_data_out[141] = ~data_out[141];
            371: correct_data_out[140] = ~data_out[140];
            372: correct_data_out[139] = ~data_out[139];
            373: correct_data_out[138] = ~data_out[138];
            374: correct_data_out[137] = ~data_out[137];
            375: correct_data_out[136] = ~data_out[136];
            376: correct_data_out[135] = ~data_out[135];
            377: correct_data_out[134] = ~data_out[134];
            378: correct_data_out[133] = ~data_out[133];
            379: correct_data_out[132] = ~data_out[132];
            380: correct_data_out[131] = ~data_out[131];
            381: correct_data_out[130] = ~data_out[130];
            382: correct_data_out[129] = ~data_out[129];
            383: correct_data_out[128] = ~data_out[128];
            384: correct_data_out[127] = ~data_out[127];
            385: correct_data_out[126] = ~data_out[126];
            386: correct_data_out[125] = ~data_out[125];
            387: correct_data_out[124] = ~data_out[124];
            388: correct_data_out[123] = ~data_out[123];
            389: correct_data_out[122] = ~data_out[122];
            390: correct_data_out[121] = ~data_out[121];
            391: correct_data_out[120] = ~data_out[120];
            392: correct_data_out[119] = ~data_out[119];
            393: correct_data_out[118] = ~data_out[118];
            394: correct_data_out[117] = ~data_out[117];
            395: correct_data_out[116] = ~data_out[116];
            396: correct_data_out[115] = ~data_out[115];
            397: correct_data_out[114] = ~data_out[114];
            398: correct_data_out[113] = ~data_out[113];
            399: correct_data_out[112] = ~data_out[112];
            400: correct_data_out[111] = ~data_out[111];
            401: correct_data_out[110] = ~data_out[110];
            402: correct_data_out[109] = ~data_out[109];
            403: correct_data_out[108] = ~data_out[108];
            404: correct_data_out[107] = ~data_out[107];
            405: correct_data_out[106] = ~data_out[106];
            406: correct_data_out[105] = ~data_out[105];
            407: correct_data_out[104] = ~data_out[104];
            408: correct_data_out[103] = ~data_out[103];
            409: correct_data_out[102] = ~data_out[102];
            410: correct_data_out[101] = ~data_out[101];
            411: correct_data_out[100] = ~data_out[100];
            412: correct_data_out[99] = ~data_out[99];
            413: correct_data_out[98] = ~data_out[98];
            414: correct_data_out[97] = ~data_out[97];
            415: correct_data_out[96] = ~data_out[96];
            416: correct_data_out[95] = ~data_out[95];
            417: correct_data_out[94] = ~data_out[94];
            418: correct_data_out[93] = ~data_out[93];
            419: correct_data_out[92] = ~data_out[92];
            420: correct_data_out[91] = ~data_out[91];
            421: correct_data_out[90] = ~data_out[90];
            422: correct_data_out[89] = ~data_out[89];
            423: correct_data_out[88] = ~data_out[88];
            424: correct_data_out[87] = ~data_out[87];
            425: correct_data_out[86] = ~data_out[86];
            426: correct_data_out[85] = ~data_out[85];
            427: correct_data_out[84] = ~data_out[84];
            428: correct_data_out[83] = ~data_out[83];
            429: correct_data_out[82] = ~data_out[82];
            430: correct_data_out[81] = ~data_out[81];
            431: correct_data_out[80] = ~data_out[80];
            432: correct_data_out[79] = ~data_out[79];
            433: correct_data_out[78] = ~data_out[78];
            434: correct_data_out[77] = ~data_out[77];
            435: correct_data_out[76] = ~data_out[76];
            436: correct_data_out[75] = ~data_out[75];
            437: correct_data_out[74] = ~data_out[74];
            438: correct_data_out[73] = ~data_out[73];
            439: correct_data_out[72] = ~data_out[72];
            440: correct_data_out[71] = ~data_out[71];
            441: correct_data_out[70] = ~data_out[70];
            442: correct_data_out[69] = ~data_out[69];
            443: correct_data_out[68] = ~data_out[68];
            444: correct_data_out[67] = ~data_out[67];
            445: correct_data_out[66] = ~data_out[66];
            446: correct_data_out[65] = ~data_out[65];
            447: correct_data_out[64] = ~data_out[64];
            448: correct_data_out[63] = ~data_out[63];
            449: correct_data_out[62] = ~data_out[62];
            450: correct_data_out[61] = ~data_out[61];
            451: correct_data_out[60] = ~data_out[60];
            452: correct_data_out[59] = ~data_out[59];
            453: correct_data_out[58] = ~data_out[58];
            454: correct_data_out[57] = ~data_out[57];
            455: correct_data_out[56] = ~data_out[56];
            456: correct_data_out[55] = ~data_out[55];
            457: correct_data_out[54] = ~data_out[54];
            458: correct_data_out[53] = ~data_out[53];
            459: correct_data_out[52] = ~data_out[52];
            460: correct_data_out[51] = ~data_out[51];
            461: correct_data_out[50] = ~data_out[50];
            462: correct_data_out[49] = ~data_out[49];
            463: correct_data_out[48] = ~data_out[48];
            464: correct_data_out[47] = ~data_out[47];
            465: correct_data_out[46] = ~data_out[46];
            466: correct_data_out[45] = ~data_out[45];
            467: correct_data_out[44] = ~data_out[44];
            468: correct_data_out[43] = ~data_out[43];
            469: correct_data_out[42] = ~data_out[42];
            470: correct_data_out[41] = ~data_out[41];
            471: correct_data_out[40] = ~data_out[40];
            472: correct_data_out[39] = ~data_out[39];
            473: correct_data_out[38] = ~data_out[38];
            474: correct_data_out[37] = ~data_out[37];
            475: correct_data_out[36] = ~data_out[36];
            476: correct_data_out[35] = ~data_out[35];
            477: correct_data_out[34] = ~data_out[34];
            478: correct_data_out[33] = ~data_out[33];
            479: correct_data_out[32] = ~data_out[32];
            480: correct_data_out[31] = ~data_out[31];
            481: correct_data_out[30] = ~data_out[30];
            482: correct_data_out[29] = ~data_out[29];
            483: correct_data_out[28] = ~data_out[28];
            484: correct_data_out[27] = ~data_out[27];
            485: correct_data_out[26] = ~data_out[26];
            486: correct_data_out[25] = ~data_out[25];
            487: correct_data_out[24] = ~data_out[24];
            488: correct_data_out[23] = ~data_out[23];
            489: correct_data_out[22] = ~data_out[22];
            490: correct_data_out[21] = ~data_out[21];
            491: correct_data_out[20] = ~data_out[20];
            492: correct_data_out[19] = ~data_out[19];
            493: correct_data_out[18] = ~data_out[18];
            494: correct_data_out[17] = ~data_out[17];
            495: correct_data_out[16] = ~data_out[16];
            496: correct_data_out[15] = ~data_out[15];
            497: correct_data_out[14] = ~data_out[14];
            498: correct_data_out[13] = ~data_out[13];
            499: correct_data_out[12] = ~data_out[12];
            500: correct_data_out[11] = ~data_out[11];
            501: correct_data_out[10] = ~data_out[10];
            502: correct_data_out[9] = ~data_out[9];
            503: correct_data_out[8] = ~data_out[8];
            504: correct_data_out[7] = ~data_out[7];
            505: correct_data_out[6] = ~data_out[6];
            506: correct_data_out[5] = ~data_out[5];
            507: correct_data_out[4] = ~data_out[4];
            508: correct_data_out[3] = ~data_out[3];
            509: correct_data_out[2] = ~data_out[2];
            510: correct_data_out[1] = ~data_out[1];
            511: correct_data_out[0] = ~data_out[0];
        endcase
    end
end // always(*)
endmodule


module mem_with_ecc_10(clock, reset, we, data_in, correct_data_out, error);

input              clock;
input              reset;
input              we;
input      [ 501:0] data_in;
output     [ 501:0] correct_data_out;
output             error;

wire       [ 501:0] data_out;
wire       [  8:0] checker_in;
wire       [  8:0] checker_out;
wire               parity_in;
wire               parity_out;

ecc_checker_10 u_checker(data_in, checker_in, parity_in);
data_mem_10 u_datamem(clock, reset, we, data_in, data_out);
ecc_mem_10 u_eccmem(clock, reset, we, checker_in, parity_in, checker_out, parity_out);
ecc_corrector_10 u_corrector(data_out, checker_out, parity_out, correct_data_out, error);

endmodule


